magic
tech sky130A
magscale 1 2
timestamp 1729373823
<< obsli1 >>
rect 1104 2159 67068 34833
<< obsm1 >>
rect 1104 552 67882 36576
<< metal2 >>
rect 4158 36551 4214 37351
rect 4342 36551 4398 37351
rect 4526 36551 4582 37351
rect 4710 36551 4766 37351
rect 4894 36551 4950 37351
rect 5078 36551 5134 37351
rect 5262 36551 5318 37351
rect 5446 36551 5502 37351
rect 5630 36551 5686 37351
rect 5814 36551 5870 37351
rect 5998 36551 6054 37351
rect 6182 36551 6238 37351
rect 6366 36551 6422 37351
rect 6550 36551 6606 37351
rect 6734 36551 6790 37351
rect 6918 36551 6974 37351
rect 7102 36551 7158 37351
rect 7286 36551 7342 37351
rect 7470 36551 7526 37351
rect 7654 36551 7710 37351
rect 7838 36551 7894 37351
rect 8022 36551 8078 37351
rect 8206 36551 8262 37351
rect 8390 36551 8446 37351
rect 8574 36551 8630 37351
rect 8758 36551 8814 37351
rect 8942 36551 8998 37351
rect 9126 36551 9182 37351
rect 9310 36551 9366 37351
rect 9494 36551 9550 37351
rect 9678 36551 9734 37351
rect 9862 36551 9918 37351
rect 10046 36551 10102 37351
rect 10230 36551 10286 37351
rect 10414 36551 10470 37351
rect 10598 36551 10654 37351
rect 10782 36551 10838 37351
rect 10966 36551 11022 37351
rect 11150 36551 11206 37351
rect 11334 36551 11390 37351
rect 11518 36551 11574 37351
rect 11702 36551 11758 37351
rect 11886 36551 11942 37351
rect 12070 36551 12126 37351
rect 12254 36551 12310 37351
rect 12438 36551 12494 37351
rect 12622 36551 12678 37351
rect 12806 36551 12862 37351
rect 12990 36551 13046 37351
rect 13174 36551 13230 37351
rect 13358 36551 13414 37351
rect 13542 36551 13598 37351
rect 13726 36551 13782 37351
rect 13910 36551 13966 37351
rect 14094 36551 14150 37351
rect 14278 36551 14334 37351
rect 14462 36551 14518 37351
rect 14646 36551 14702 37351
rect 14830 36551 14886 37351
rect 15014 36551 15070 37351
rect 15198 36551 15254 37351
rect 15382 36551 15438 37351
rect 15566 36551 15622 37351
rect 15750 36551 15806 37351
rect 15934 36551 15990 37351
rect 16118 36551 16174 37351
rect 16302 36551 16358 37351
rect 16486 36551 16542 37351
rect 16670 36551 16726 37351
rect 16854 36551 16910 37351
rect 17038 36551 17094 37351
rect 17222 36551 17278 37351
rect 17406 36551 17462 37351
rect 17590 36551 17646 37351
rect 17774 36551 17830 37351
rect 17958 36551 18014 37351
rect 18142 36551 18198 37351
rect 18326 36551 18382 37351
rect 18510 36551 18566 37351
rect 18694 36551 18750 37351
rect 18878 36551 18934 37351
rect 19062 36551 19118 37351
rect 19246 36551 19302 37351
rect 19430 36551 19486 37351
rect 19614 36551 19670 37351
rect 19798 36551 19854 37351
rect 19982 36551 20038 37351
rect 20166 36551 20222 37351
rect 20350 36551 20406 37351
rect 20534 36551 20590 37351
rect 20718 36551 20774 37351
rect 20902 36551 20958 37351
rect 21086 36551 21142 37351
rect 21270 36551 21326 37351
rect 21454 36551 21510 37351
rect 21638 36551 21694 37351
rect 21822 36551 21878 37351
rect 22006 36551 22062 37351
rect 22190 36551 22246 37351
rect 22374 36551 22430 37351
rect 22558 36551 22614 37351
rect 22742 36551 22798 37351
rect 22926 36551 22982 37351
rect 23110 36551 23166 37351
rect 23294 36551 23350 37351
rect 23478 36551 23534 37351
rect 23662 36551 23718 37351
rect 23846 36551 23902 37351
rect 24030 36551 24086 37351
rect 24214 36551 24270 37351
rect 24398 36551 24454 37351
rect 24582 36551 24638 37351
rect 24766 36551 24822 37351
rect 24950 36551 25006 37351
rect 25134 36551 25190 37351
rect 25318 36551 25374 37351
rect 25502 36551 25558 37351
rect 25686 36551 25742 37351
rect 25870 36551 25926 37351
rect 26054 36551 26110 37351
rect 26238 36551 26294 37351
rect 26422 36551 26478 37351
rect 26606 36551 26662 37351
rect 26790 36551 26846 37351
rect 26974 36551 27030 37351
rect 27158 36551 27214 37351
rect 27342 36551 27398 37351
rect 27526 36551 27582 37351
rect 27710 36551 27766 37351
rect 27894 36551 27950 37351
rect 28078 36551 28134 37351
rect 28262 36551 28318 37351
rect 28446 36551 28502 37351
rect 28630 36551 28686 37351
rect 28814 36551 28870 37351
rect 28998 36551 29054 37351
rect 29182 36551 29238 37351
rect 29366 36551 29422 37351
rect 29550 36551 29606 37351
rect 29734 36551 29790 37351
rect 29918 36551 29974 37351
rect 30102 36551 30158 37351
rect 30286 36551 30342 37351
rect 30470 36551 30526 37351
rect 30654 36551 30710 37351
rect 30838 36551 30894 37351
rect 31022 36551 31078 37351
rect 31206 36551 31262 37351
rect 31390 36551 31446 37351
rect 31574 36551 31630 37351
rect 31758 36551 31814 37351
rect 31942 36551 31998 37351
rect 32126 36551 32182 37351
rect 32310 36551 32366 37351
rect 32494 36551 32550 37351
rect 32678 36551 32734 37351
rect 32862 36551 32918 37351
rect 33046 36551 33102 37351
rect 33230 36551 33286 37351
rect 33414 36551 33470 37351
rect 33598 36551 33654 37351
rect 33782 36551 33838 37351
rect 33966 36551 34022 37351
rect 34150 36551 34206 37351
rect 34334 36551 34390 37351
rect 34518 36551 34574 37351
rect 34702 36551 34758 37351
rect 34886 36551 34942 37351
rect 35070 36551 35126 37351
rect 35254 36551 35310 37351
rect 35438 36551 35494 37351
rect 35622 36551 35678 37351
rect 35806 36551 35862 37351
rect 35990 36551 36046 37351
rect 36174 36551 36230 37351
rect 36358 36551 36414 37351
rect 36542 36551 36598 37351
rect 36726 36551 36782 37351
rect 36910 36551 36966 37351
rect 37094 36551 37150 37351
rect 37278 36551 37334 37351
rect 37462 36551 37518 37351
rect 37646 36551 37702 37351
rect 37830 36551 37886 37351
rect 38014 36551 38070 37351
rect 38198 36551 38254 37351
rect 38382 36551 38438 37351
rect 38566 36551 38622 37351
rect 38750 36551 38806 37351
rect 38934 36551 38990 37351
rect 39118 36551 39174 37351
rect 39302 36551 39358 37351
rect 39486 36551 39542 37351
rect 39670 36551 39726 37351
rect 39854 36551 39910 37351
rect 40038 36551 40094 37351
rect 40222 36551 40278 37351
rect 40406 36551 40462 37351
rect 40590 36551 40646 37351
rect 40774 36551 40830 37351
rect 40958 36551 41014 37351
rect 41142 36551 41198 37351
rect 41326 36551 41382 37351
rect 41510 36551 41566 37351
rect 41694 36551 41750 37351
rect 41878 36551 41934 37351
rect 42062 36551 42118 37351
rect 42246 36551 42302 37351
rect 42430 36551 42486 37351
rect 42614 36551 42670 37351
rect 42798 36551 42854 37351
rect 42982 36551 43038 37351
rect 43166 36551 43222 37351
rect 43350 36551 43406 37351
rect 43534 36551 43590 37351
rect 43718 36551 43774 37351
rect 43902 36551 43958 37351
rect 44086 36551 44142 37351
rect 44270 36551 44326 37351
rect 44454 36551 44510 37351
rect 44638 36551 44694 37351
rect 44822 36551 44878 37351
rect 45006 36551 45062 37351
rect 45190 36551 45246 37351
rect 45374 36551 45430 37351
rect 45558 36551 45614 37351
rect 45742 36551 45798 37351
rect 45926 36551 45982 37351
rect 46110 36551 46166 37351
rect 46294 36551 46350 37351
rect 46478 36551 46534 37351
rect 46662 36551 46718 37351
rect 46846 36551 46902 37351
rect 47030 36551 47086 37351
rect 47214 36551 47270 37351
rect 47398 36551 47454 37351
rect 47582 36551 47638 37351
rect 47766 36551 47822 37351
rect 47950 36551 48006 37351
rect 48134 36551 48190 37351
rect 48318 36551 48374 37351
rect 48502 36551 48558 37351
rect 48686 36551 48742 37351
rect 48870 36551 48926 37351
rect 49054 36551 49110 37351
rect 49238 36551 49294 37351
rect 49422 36551 49478 37351
rect 49606 36551 49662 37351
rect 49790 36551 49846 37351
rect 49974 36551 50030 37351
rect 50158 36551 50214 37351
rect 50342 36551 50398 37351
rect 50526 36551 50582 37351
rect 50710 36551 50766 37351
rect 50894 36551 50950 37351
rect 51078 36551 51134 37351
rect 51262 36551 51318 37351
rect 51446 36551 51502 37351
rect 51630 36551 51686 37351
rect 51814 36551 51870 37351
rect 51998 36551 52054 37351
rect 52182 36551 52238 37351
rect 52366 36551 52422 37351
rect 52550 36551 52606 37351
rect 52734 36551 52790 37351
rect 52918 36551 52974 37351
rect 53102 36551 53158 37351
rect 53286 36551 53342 37351
rect 53470 36551 53526 37351
rect 53654 36551 53710 37351
rect 53838 36551 53894 37351
rect 54022 36551 54078 37351
rect 54206 36551 54262 37351
rect 54390 36551 54446 37351
rect 54574 36551 54630 37351
rect 54758 36551 54814 37351
rect 54942 36551 54998 37351
rect 55126 36551 55182 37351
rect 55310 36551 55366 37351
rect 55494 36551 55550 37351
rect 55678 36551 55734 37351
rect 55862 36551 55918 37351
rect 56046 36551 56102 37351
rect 56230 36551 56286 37351
rect 56414 36551 56470 37351
rect 56598 36551 56654 37351
rect 56782 36551 56838 37351
rect 56966 36551 57022 37351
rect 57150 36551 57206 37351
rect 57334 36551 57390 37351
rect 57518 36551 57574 37351
rect 57702 36551 57758 37351
rect 57886 36551 57942 37351
rect 58070 36551 58126 37351
rect 58254 36551 58310 37351
rect 58438 36551 58494 37351
rect 58622 36551 58678 37351
rect 58806 36551 58862 37351
rect 58990 36551 59046 37351
rect 59174 36551 59230 37351
rect 59358 36551 59414 37351
rect 59542 36551 59598 37351
rect 59726 36551 59782 37351
rect 59910 36551 59966 37351
rect 60094 36551 60150 37351
rect 60278 36551 60334 37351
rect 60462 36551 60518 37351
rect 60646 36551 60702 37351
rect 60830 36551 60886 37351
rect 61014 36551 61070 37351
rect 61198 36551 61254 37351
rect 61382 36551 61438 37351
rect 61566 36551 61622 37351
rect 61750 36551 61806 37351
rect 61934 36551 61990 37351
rect 62118 36551 62174 37351
rect 62302 36551 62358 37351
rect 62486 36551 62542 37351
rect 62670 36551 62726 37351
rect 62854 36551 62910 37351
rect 63038 36551 63094 37351
rect 63222 36551 63278 37351
rect 63406 36551 63462 37351
rect 63590 36551 63646 37351
rect 63774 36551 63830 37351
rect 63958 36551 64014 37351
rect 10414 0 10470 800
rect 10598 0 10654 800
rect 10782 0 10838 800
rect 10966 0 11022 800
rect 11150 0 11206 800
rect 11334 0 11390 800
rect 11518 0 11574 800
rect 11702 0 11758 800
rect 11886 0 11942 800
rect 12070 0 12126 800
rect 12254 0 12310 800
rect 12438 0 12494 800
rect 12622 0 12678 800
rect 12806 0 12862 800
rect 12990 0 13046 800
rect 13174 0 13230 800
rect 13358 0 13414 800
rect 13542 0 13598 800
rect 13726 0 13782 800
rect 13910 0 13966 800
rect 14094 0 14150 800
rect 14278 0 14334 800
rect 14462 0 14518 800
rect 14646 0 14702 800
rect 14830 0 14886 800
rect 15014 0 15070 800
rect 15198 0 15254 800
rect 15382 0 15438 800
rect 15566 0 15622 800
rect 15750 0 15806 800
rect 15934 0 15990 800
rect 16118 0 16174 800
rect 16302 0 16358 800
rect 16486 0 16542 800
rect 16670 0 16726 800
rect 16854 0 16910 800
rect 17038 0 17094 800
rect 17222 0 17278 800
rect 17406 0 17462 800
rect 17590 0 17646 800
rect 17774 0 17830 800
rect 17958 0 18014 800
rect 18142 0 18198 800
rect 18326 0 18382 800
rect 18510 0 18566 800
rect 18694 0 18750 800
rect 18878 0 18934 800
rect 19062 0 19118 800
rect 19246 0 19302 800
rect 19430 0 19486 800
rect 19614 0 19670 800
rect 19798 0 19854 800
rect 19982 0 20038 800
rect 20166 0 20222 800
rect 20350 0 20406 800
rect 20534 0 20590 800
rect 20718 0 20774 800
rect 20902 0 20958 800
rect 21086 0 21142 800
rect 21270 0 21326 800
rect 21454 0 21510 800
rect 21638 0 21694 800
rect 21822 0 21878 800
rect 22006 0 22062 800
rect 22190 0 22246 800
rect 22374 0 22430 800
rect 22558 0 22614 800
rect 22742 0 22798 800
rect 22926 0 22982 800
rect 23110 0 23166 800
rect 23294 0 23350 800
rect 23478 0 23534 800
rect 23662 0 23718 800
rect 23846 0 23902 800
rect 24030 0 24086 800
rect 24214 0 24270 800
rect 24398 0 24454 800
rect 24582 0 24638 800
rect 24766 0 24822 800
rect 24950 0 25006 800
rect 25134 0 25190 800
rect 25318 0 25374 800
rect 25502 0 25558 800
rect 25686 0 25742 800
rect 25870 0 25926 800
rect 26054 0 26110 800
rect 26238 0 26294 800
rect 26422 0 26478 800
rect 26606 0 26662 800
rect 26790 0 26846 800
rect 26974 0 27030 800
rect 27158 0 27214 800
rect 27342 0 27398 800
rect 27526 0 27582 800
rect 27710 0 27766 800
rect 27894 0 27950 800
rect 28078 0 28134 800
rect 28262 0 28318 800
rect 28446 0 28502 800
rect 28630 0 28686 800
rect 28814 0 28870 800
rect 28998 0 29054 800
rect 29182 0 29238 800
rect 29366 0 29422 800
rect 29550 0 29606 800
rect 29734 0 29790 800
rect 29918 0 29974 800
rect 30102 0 30158 800
rect 30286 0 30342 800
rect 30470 0 30526 800
rect 30654 0 30710 800
rect 30838 0 30894 800
rect 31022 0 31078 800
rect 31206 0 31262 800
rect 31390 0 31446 800
rect 31574 0 31630 800
rect 31758 0 31814 800
rect 31942 0 31998 800
rect 32126 0 32182 800
rect 32310 0 32366 800
rect 32494 0 32550 800
rect 32678 0 32734 800
rect 32862 0 32918 800
rect 33046 0 33102 800
rect 33230 0 33286 800
rect 33414 0 33470 800
rect 33598 0 33654 800
rect 33782 0 33838 800
rect 33966 0 34022 800
rect 34150 0 34206 800
rect 34334 0 34390 800
rect 34518 0 34574 800
rect 34702 0 34758 800
rect 34886 0 34942 800
rect 35070 0 35126 800
rect 35254 0 35310 800
rect 35438 0 35494 800
rect 35622 0 35678 800
rect 35806 0 35862 800
rect 35990 0 36046 800
rect 36174 0 36230 800
rect 36358 0 36414 800
rect 36542 0 36598 800
rect 36726 0 36782 800
rect 36910 0 36966 800
rect 37094 0 37150 800
rect 37278 0 37334 800
rect 37462 0 37518 800
rect 37646 0 37702 800
rect 37830 0 37886 800
rect 38014 0 38070 800
rect 38198 0 38254 800
rect 38382 0 38438 800
rect 38566 0 38622 800
rect 38750 0 38806 800
rect 38934 0 38990 800
rect 39118 0 39174 800
rect 39302 0 39358 800
rect 39486 0 39542 800
rect 39670 0 39726 800
rect 39854 0 39910 800
rect 40038 0 40094 800
rect 40222 0 40278 800
rect 40406 0 40462 800
rect 40590 0 40646 800
rect 40774 0 40830 800
rect 40958 0 41014 800
rect 41142 0 41198 800
rect 41326 0 41382 800
rect 41510 0 41566 800
rect 41694 0 41750 800
rect 41878 0 41934 800
rect 42062 0 42118 800
rect 42246 0 42302 800
rect 42430 0 42486 800
rect 42614 0 42670 800
rect 42798 0 42854 800
rect 42982 0 43038 800
rect 43166 0 43222 800
rect 43350 0 43406 800
rect 43534 0 43590 800
rect 43718 0 43774 800
rect 43902 0 43958 800
rect 44086 0 44142 800
rect 44270 0 44326 800
rect 44454 0 44510 800
rect 44638 0 44694 800
rect 44822 0 44878 800
rect 45006 0 45062 800
rect 45190 0 45246 800
rect 45374 0 45430 800
rect 45558 0 45614 800
rect 45742 0 45798 800
rect 45926 0 45982 800
rect 46110 0 46166 800
rect 46294 0 46350 800
rect 46478 0 46534 800
rect 46662 0 46718 800
rect 46846 0 46902 800
rect 47030 0 47086 800
rect 47214 0 47270 800
rect 47398 0 47454 800
rect 47582 0 47638 800
rect 47766 0 47822 800
rect 47950 0 48006 800
rect 48134 0 48190 800
rect 48318 0 48374 800
rect 48502 0 48558 800
rect 48686 0 48742 800
rect 48870 0 48926 800
rect 49054 0 49110 800
rect 49238 0 49294 800
rect 49422 0 49478 800
rect 49606 0 49662 800
rect 49790 0 49846 800
rect 49974 0 50030 800
rect 50158 0 50214 800
rect 50342 0 50398 800
rect 50526 0 50582 800
rect 50710 0 50766 800
rect 50894 0 50950 800
rect 51078 0 51134 800
rect 51262 0 51318 800
rect 51446 0 51502 800
rect 51630 0 51686 800
rect 51814 0 51870 800
rect 51998 0 52054 800
rect 52182 0 52238 800
rect 52366 0 52422 800
rect 52550 0 52606 800
rect 52734 0 52790 800
rect 52918 0 52974 800
rect 53102 0 53158 800
rect 53286 0 53342 800
rect 53470 0 53526 800
rect 53654 0 53710 800
rect 53838 0 53894 800
rect 54022 0 54078 800
rect 54206 0 54262 800
rect 54390 0 54446 800
rect 54574 0 54630 800
rect 54758 0 54814 800
rect 54942 0 54998 800
rect 55126 0 55182 800
rect 55310 0 55366 800
rect 55494 0 55550 800
rect 55678 0 55734 800
rect 55862 0 55918 800
rect 56046 0 56102 800
rect 56230 0 56286 800
rect 56414 0 56470 800
rect 56598 0 56654 800
rect 56782 0 56838 800
rect 56966 0 57022 800
rect 57150 0 57206 800
rect 57334 0 57390 800
rect 57518 0 57574 800
rect 57702 0 57758 800
<< obsm2 >>
rect 1214 36495 4102 36666
rect 4270 36495 4286 36666
rect 4454 36495 4470 36666
rect 4638 36495 4654 36666
rect 4822 36495 4838 36666
rect 5006 36495 5022 36666
rect 5190 36495 5206 36666
rect 5374 36495 5390 36666
rect 5558 36495 5574 36666
rect 5742 36495 5758 36666
rect 5926 36495 5942 36666
rect 6110 36495 6126 36666
rect 6294 36495 6310 36666
rect 6478 36495 6494 36666
rect 6662 36495 6678 36666
rect 6846 36495 6862 36666
rect 7030 36495 7046 36666
rect 7214 36495 7230 36666
rect 7398 36495 7414 36666
rect 7582 36495 7598 36666
rect 7766 36495 7782 36666
rect 7950 36495 7966 36666
rect 8134 36495 8150 36666
rect 8318 36495 8334 36666
rect 8502 36495 8518 36666
rect 8686 36495 8702 36666
rect 8870 36495 8886 36666
rect 9054 36495 9070 36666
rect 9238 36495 9254 36666
rect 9422 36495 9438 36666
rect 9606 36495 9622 36666
rect 9790 36495 9806 36666
rect 9974 36495 9990 36666
rect 10158 36495 10174 36666
rect 10342 36495 10358 36666
rect 10526 36495 10542 36666
rect 10710 36495 10726 36666
rect 10894 36495 10910 36666
rect 11078 36495 11094 36666
rect 11262 36495 11278 36666
rect 11446 36495 11462 36666
rect 11630 36495 11646 36666
rect 11814 36495 11830 36666
rect 11998 36495 12014 36666
rect 12182 36495 12198 36666
rect 12366 36495 12382 36666
rect 12550 36495 12566 36666
rect 12734 36495 12750 36666
rect 12918 36495 12934 36666
rect 13102 36495 13118 36666
rect 13286 36495 13302 36666
rect 13470 36495 13486 36666
rect 13654 36495 13670 36666
rect 13838 36495 13854 36666
rect 14022 36495 14038 36666
rect 14206 36495 14222 36666
rect 14390 36495 14406 36666
rect 14574 36495 14590 36666
rect 14758 36495 14774 36666
rect 14942 36495 14958 36666
rect 15126 36495 15142 36666
rect 15310 36495 15326 36666
rect 15494 36495 15510 36666
rect 15678 36495 15694 36666
rect 15862 36495 15878 36666
rect 16046 36495 16062 36666
rect 16230 36495 16246 36666
rect 16414 36495 16430 36666
rect 16598 36495 16614 36666
rect 16782 36495 16798 36666
rect 16966 36495 16982 36666
rect 17150 36495 17166 36666
rect 17334 36495 17350 36666
rect 17518 36495 17534 36666
rect 17702 36495 17718 36666
rect 17886 36495 17902 36666
rect 18070 36495 18086 36666
rect 18254 36495 18270 36666
rect 18438 36495 18454 36666
rect 18622 36495 18638 36666
rect 18806 36495 18822 36666
rect 18990 36495 19006 36666
rect 19174 36495 19190 36666
rect 19358 36495 19374 36666
rect 19542 36495 19558 36666
rect 19726 36495 19742 36666
rect 19910 36495 19926 36666
rect 20094 36495 20110 36666
rect 20278 36495 20294 36666
rect 20462 36495 20478 36666
rect 20646 36495 20662 36666
rect 20830 36495 20846 36666
rect 21014 36495 21030 36666
rect 21198 36495 21214 36666
rect 21382 36495 21398 36666
rect 21566 36495 21582 36666
rect 21750 36495 21766 36666
rect 21934 36495 21950 36666
rect 22118 36495 22134 36666
rect 22302 36495 22318 36666
rect 22486 36495 22502 36666
rect 22670 36495 22686 36666
rect 22854 36495 22870 36666
rect 23038 36495 23054 36666
rect 23222 36495 23238 36666
rect 23406 36495 23422 36666
rect 23590 36495 23606 36666
rect 23774 36495 23790 36666
rect 23958 36495 23974 36666
rect 24142 36495 24158 36666
rect 24326 36495 24342 36666
rect 24510 36495 24526 36666
rect 24694 36495 24710 36666
rect 24878 36495 24894 36666
rect 25062 36495 25078 36666
rect 25246 36495 25262 36666
rect 25430 36495 25446 36666
rect 25614 36495 25630 36666
rect 25798 36495 25814 36666
rect 25982 36495 25998 36666
rect 26166 36495 26182 36666
rect 26350 36495 26366 36666
rect 26534 36495 26550 36666
rect 26718 36495 26734 36666
rect 26902 36495 26918 36666
rect 27086 36495 27102 36666
rect 27270 36495 27286 36666
rect 27454 36495 27470 36666
rect 27638 36495 27654 36666
rect 27822 36495 27838 36666
rect 28006 36495 28022 36666
rect 28190 36495 28206 36666
rect 28374 36495 28390 36666
rect 28558 36495 28574 36666
rect 28742 36495 28758 36666
rect 28926 36495 28942 36666
rect 29110 36495 29126 36666
rect 29294 36495 29310 36666
rect 29478 36495 29494 36666
rect 29662 36495 29678 36666
rect 29846 36495 29862 36666
rect 30030 36495 30046 36666
rect 30214 36495 30230 36666
rect 30398 36495 30414 36666
rect 30582 36495 30598 36666
rect 30766 36495 30782 36666
rect 30950 36495 30966 36666
rect 31134 36495 31150 36666
rect 31318 36495 31334 36666
rect 31502 36495 31518 36666
rect 31686 36495 31702 36666
rect 31870 36495 31886 36666
rect 32054 36495 32070 36666
rect 32238 36495 32254 36666
rect 32422 36495 32438 36666
rect 32606 36495 32622 36666
rect 32790 36495 32806 36666
rect 32974 36495 32990 36666
rect 33158 36495 33174 36666
rect 33342 36495 33358 36666
rect 33526 36495 33542 36666
rect 33710 36495 33726 36666
rect 33894 36495 33910 36666
rect 34078 36495 34094 36666
rect 34262 36495 34278 36666
rect 34446 36495 34462 36666
rect 34630 36495 34646 36666
rect 34814 36495 34830 36666
rect 34998 36495 35014 36666
rect 35182 36495 35198 36666
rect 35366 36495 35382 36666
rect 35550 36495 35566 36666
rect 35734 36495 35750 36666
rect 35918 36495 35934 36666
rect 36102 36495 36118 36666
rect 36286 36495 36302 36666
rect 36470 36495 36486 36666
rect 36654 36495 36670 36666
rect 36838 36495 36854 36666
rect 37022 36495 37038 36666
rect 37206 36495 37222 36666
rect 37390 36495 37406 36666
rect 37574 36495 37590 36666
rect 37758 36495 37774 36666
rect 37942 36495 37958 36666
rect 38126 36495 38142 36666
rect 38310 36495 38326 36666
rect 38494 36495 38510 36666
rect 38678 36495 38694 36666
rect 38862 36495 38878 36666
rect 39046 36495 39062 36666
rect 39230 36495 39246 36666
rect 39414 36495 39430 36666
rect 39598 36495 39614 36666
rect 39782 36495 39798 36666
rect 39966 36495 39982 36666
rect 40150 36495 40166 36666
rect 40334 36495 40350 36666
rect 40518 36495 40534 36666
rect 40702 36495 40718 36666
rect 40886 36495 40902 36666
rect 41070 36495 41086 36666
rect 41254 36495 41270 36666
rect 41438 36495 41454 36666
rect 41622 36495 41638 36666
rect 41806 36495 41822 36666
rect 41990 36495 42006 36666
rect 42174 36495 42190 36666
rect 42358 36495 42374 36666
rect 42542 36495 42558 36666
rect 42726 36495 42742 36666
rect 42910 36495 42926 36666
rect 43094 36495 43110 36666
rect 43278 36495 43294 36666
rect 43462 36495 43478 36666
rect 43646 36495 43662 36666
rect 43830 36495 43846 36666
rect 44014 36495 44030 36666
rect 44198 36495 44214 36666
rect 44382 36495 44398 36666
rect 44566 36495 44582 36666
rect 44750 36495 44766 36666
rect 44934 36495 44950 36666
rect 45118 36495 45134 36666
rect 45302 36495 45318 36666
rect 45486 36495 45502 36666
rect 45670 36495 45686 36666
rect 45854 36495 45870 36666
rect 46038 36495 46054 36666
rect 46222 36495 46238 36666
rect 46406 36495 46422 36666
rect 46590 36495 46606 36666
rect 46774 36495 46790 36666
rect 46958 36495 46974 36666
rect 47142 36495 47158 36666
rect 47326 36495 47342 36666
rect 47510 36495 47526 36666
rect 47694 36495 47710 36666
rect 47878 36495 47894 36666
rect 48062 36495 48078 36666
rect 48246 36495 48262 36666
rect 48430 36495 48446 36666
rect 48614 36495 48630 36666
rect 48798 36495 48814 36666
rect 48982 36495 48998 36666
rect 49166 36495 49182 36666
rect 49350 36495 49366 36666
rect 49534 36495 49550 36666
rect 49718 36495 49734 36666
rect 49902 36495 49918 36666
rect 50086 36495 50102 36666
rect 50270 36495 50286 36666
rect 50454 36495 50470 36666
rect 50638 36495 50654 36666
rect 50822 36495 50838 36666
rect 51006 36495 51022 36666
rect 51190 36495 51206 36666
rect 51374 36495 51390 36666
rect 51558 36495 51574 36666
rect 51742 36495 51758 36666
rect 51926 36495 51942 36666
rect 52110 36495 52126 36666
rect 52294 36495 52310 36666
rect 52478 36495 52494 36666
rect 52662 36495 52678 36666
rect 52846 36495 52862 36666
rect 53030 36495 53046 36666
rect 53214 36495 53230 36666
rect 53398 36495 53414 36666
rect 53582 36495 53598 36666
rect 53766 36495 53782 36666
rect 53950 36495 53966 36666
rect 54134 36495 54150 36666
rect 54318 36495 54334 36666
rect 54502 36495 54518 36666
rect 54686 36495 54702 36666
rect 54870 36495 54886 36666
rect 55054 36495 55070 36666
rect 55238 36495 55254 36666
rect 55422 36495 55438 36666
rect 55606 36495 55622 36666
rect 55790 36495 55806 36666
rect 55974 36495 55990 36666
rect 56158 36495 56174 36666
rect 56342 36495 56358 36666
rect 56526 36495 56542 36666
rect 56710 36495 56726 36666
rect 56894 36495 56910 36666
rect 57078 36495 57094 36666
rect 57262 36495 57278 36666
rect 57446 36495 57462 36666
rect 57630 36495 57646 36666
rect 57814 36495 57830 36666
rect 57998 36495 58014 36666
rect 58182 36495 58198 36666
rect 58366 36495 58382 36666
rect 58550 36495 58566 36666
rect 58734 36495 58750 36666
rect 58918 36495 58934 36666
rect 59102 36495 59118 36666
rect 59286 36495 59302 36666
rect 59470 36495 59486 36666
rect 59654 36495 59670 36666
rect 59838 36495 59854 36666
rect 60022 36495 60038 36666
rect 60206 36495 60222 36666
rect 60390 36495 60406 36666
rect 60574 36495 60590 36666
rect 60758 36495 60774 36666
rect 60942 36495 60958 36666
rect 61126 36495 61142 36666
rect 61310 36495 61326 36666
rect 61494 36495 61510 36666
rect 61678 36495 61694 36666
rect 61862 36495 61878 36666
rect 62046 36495 62062 36666
rect 62230 36495 62246 36666
rect 62414 36495 62430 36666
rect 62598 36495 62614 36666
rect 62782 36495 62798 36666
rect 62966 36495 62982 36666
rect 63150 36495 63166 36666
rect 63334 36495 63350 36666
rect 63518 36495 63534 36666
rect 63702 36495 63718 36666
rect 63886 36495 63902 36666
rect 64070 36495 67876 36666
rect 1214 856 67876 36495
rect 1214 546 10358 856
rect 10526 546 10542 856
rect 10710 546 10726 856
rect 10894 546 10910 856
rect 11078 546 11094 856
rect 11262 546 11278 856
rect 11446 546 11462 856
rect 11630 546 11646 856
rect 11814 546 11830 856
rect 11998 546 12014 856
rect 12182 546 12198 856
rect 12366 546 12382 856
rect 12550 546 12566 856
rect 12734 546 12750 856
rect 12918 546 12934 856
rect 13102 546 13118 856
rect 13286 546 13302 856
rect 13470 546 13486 856
rect 13654 546 13670 856
rect 13838 546 13854 856
rect 14022 546 14038 856
rect 14206 546 14222 856
rect 14390 546 14406 856
rect 14574 546 14590 856
rect 14758 546 14774 856
rect 14942 546 14958 856
rect 15126 546 15142 856
rect 15310 546 15326 856
rect 15494 546 15510 856
rect 15678 546 15694 856
rect 15862 546 15878 856
rect 16046 546 16062 856
rect 16230 546 16246 856
rect 16414 546 16430 856
rect 16598 546 16614 856
rect 16782 546 16798 856
rect 16966 546 16982 856
rect 17150 546 17166 856
rect 17334 546 17350 856
rect 17518 546 17534 856
rect 17702 546 17718 856
rect 17886 546 17902 856
rect 18070 546 18086 856
rect 18254 546 18270 856
rect 18438 546 18454 856
rect 18622 546 18638 856
rect 18806 546 18822 856
rect 18990 546 19006 856
rect 19174 546 19190 856
rect 19358 546 19374 856
rect 19542 546 19558 856
rect 19726 546 19742 856
rect 19910 546 19926 856
rect 20094 546 20110 856
rect 20278 546 20294 856
rect 20462 546 20478 856
rect 20646 546 20662 856
rect 20830 546 20846 856
rect 21014 546 21030 856
rect 21198 546 21214 856
rect 21382 546 21398 856
rect 21566 546 21582 856
rect 21750 546 21766 856
rect 21934 546 21950 856
rect 22118 546 22134 856
rect 22302 546 22318 856
rect 22486 546 22502 856
rect 22670 546 22686 856
rect 22854 546 22870 856
rect 23038 546 23054 856
rect 23222 546 23238 856
rect 23406 546 23422 856
rect 23590 546 23606 856
rect 23774 546 23790 856
rect 23958 546 23974 856
rect 24142 546 24158 856
rect 24326 546 24342 856
rect 24510 546 24526 856
rect 24694 546 24710 856
rect 24878 546 24894 856
rect 25062 546 25078 856
rect 25246 546 25262 856
rect 25430 546 25446 856
rect 25614 546 25630 856
rect 25798 546 25814 856
rect 25982 546 25998 856
rect 26166 546 26182 856
rect 26350 546 26366 856
rect 26534 546 26550 856
rect 26718 546 26734 856
rect 26902 546 26918 856
rect 27086 546 27102 856
rect 27270 546 27286 856
rect 27454 546 27470 856
rect 27638 546 27654 856
rect 27822 546 27838 856
rect 28006 546 28022 856
rect 28190 546 28206 856
rect 28374 546 28390 856
rect 28558 546 28574 856
rect 28742 546 28758 856
rect 28926 546 28942 856
rect 29110 546 29126 856
rect 29294 546 29310 856
rect 29478 546 29494 856
rect 29662 546 29678 856
rect 29846 546 29862 856
rect 30030 546 30046 856
rect 30214 546 30230 856
rect 30398 546 30414 856
rect 30582 546 30598 856
rect 30766 546 30782 856
rect 30950 546 30966 856
rect 31134 546 31150 856
rect 31318 546 31334 856
rect 31502 546 31518 856
rect 31686 546 31702 856
rect 31870 546 31886 856
rect 32054 546 32070 856
rect 32238 546 32254 856
rect 32422 546 32438 856
rect 32606 546 32622 856
rect 32790 546 32806 856
rect 32974 546 32990 856
rect 33158 546 33174 856
rect 33342 546 33358 856
rect 33526 546 33542 856
rect 33710 546 33726 856
rect 33894 546 33910 856
rect 34078 546 34094 856
rect 34262 546 34278 856
rect 34446 546 34462 856
rect 34630 546 34646 856
rect 34814 546 34830 856
rect 34998 546 35014 856
rect 35182 546 35198 856
rect 35366 546 35382 856
rect 35550 546 35566 856
rect 35734 546 35750 856
rect 35918 546 35934 856
rect 36102 546 36118 856
rect 36286 546 36302 856
rect 36470 546 36486 856
rect 36654 546 36670 856
rect 36838 546 36854 856
rect 37022 546 37038 856
rect 37206 546 37222 856
rect 37390 546 37406 856
rect 37574 546 37590 856
rect 37758 546 37774 856
rect 37942 546 37958 856
rect 38126 546 38142 856
rect 38310 546 38326 856
rect 38494 546 38510 856
rect 38678 546 38694 856
rect 38862 546 38878 856
rect 39046 546 39062 856
rect 39230 546 39246 856
rect 39414 546 39430 856
rect 39598 546 39614 856
rect 39782 546 39798 856
rect 39966 546 39982 856
rect 40150 546 40166 856
rect 40334 546 40350 856
rect 40518 546 40534 856
rect 40702 546 40718 856
rect 40886 546 40902 856
rect 41070 546 41086 856
rect 41254 546 41270 856
rect 41438 546 41454 856
rect 41622 546 41638 856
rect 41806 546 41822 856
rect 41990 546 42006 856
rect 42174 546 42190 856
rect 42358 546 42374 856
rect 42542 546 42558 856
rect 42726 546 42742 856
rect 42910 546 42926 856
rect 43094 546 43110 856
rect 43278 546 43294 856
rect 43462 546 43478 856
rect 43646 546 43662 856
rect 43830 546 43846 856
rect 44014 546 44030 856
rect 44198 546 44214 856
rect 44382 546 44398 856
rect 44566 546 44582 856
rect 44750 546 44766 856
rect 44934 546 44950 856
rect 45118 546 45134 856
rect 45302 546 45318 856
rect 45486 546 45502 856
rect 45670 546 45686 856
rect 45854 546 45870 856
rect 46038 546 46054 856
rect 46222 546 46238 856
rect 46406 546 46422 856
rect 46590 546 46606 856
rect 46774 546 46790 856
rect 46958 546 46974 856
rect 47142 546 47158 856
rect 47326 546 47342 856
rect 47510 546 47526 856
rect 47694 546 47710 856
rect 47878 546 47894 856
rect 48062 546 48078 856
rect 48246 546 48262 856
rect 48430 546 48446 856
rect 48614 546 48630 856
rect 48798 546 48814 856
rect 48982 546 48998 856
rect 49166 546 49182 856
rect 49350 546 49366 856
rect 49534 546 49550 856
rect 49718 546 49734 856
rect 49902 546 49918 856
rect 50086 546 50102 856
rect 50270 546 50286 856
rect 50454 546 50470 856
rect 50638 546 50654 856
rect 50822 546 50838 856
rect 51006 546 51022 856
rect 51190 546 51206 856
rect 51374 546 51390 856
rect 51558 546 51574 856
rect 51742 546 51758 856
rect 51926 546 51942 856
rect 52110 546 52126 856
rect 52294 546 52310 856
rect 52478 546 52494 856
rect 52662 546 52678 856
rect 52846 546 52862 856
rect 53030 546 53046 856
rect 53214 546 53230 856
rect 53398 546 53414 856
rect 53582 546 53598 856
rect 53766 546 53782 856
rect 53950 546 53966 856
rect 54134 546 54150 856
rect 54318 546 54334 856
rect 54502 546 54518 856
rect 54686 546 54702 856
rect 54870 546 54886 856
rect 55054 546 55070 856
rect 55238 546 55254 856
rect 55422 546 55438 856
rect 55606 546 55622 856
rect 55790 546 55806 856
rect 55974 546 55990 856
rect 56158 546 56174 856
rect 56342 546 56358 856
rect 56526 546 56542 856
rect 56710 546 56726 856
rect 56894 546 56910 856
rect 57078 546 57094 856
rect 57262 546 57278 856
rect 57446 546 57462 856
rect 57630 546 57646 856
rect 57814 546 67876 856
<< metal3 >>
rect 0 36184 800 36304
rect 0 35640 800 35760
rect 0 35096 800 35216
rect 0 34552 800 34672
rect 0 34008 800 34128
rect 0 33464 800 33584
rect 0 32920 800 33040
rect 0 32376 800 32496
rect 0 31832 800 31952
rect 0 31288 800 31408
rect 0 30744 800 30864
rect 0 30200 800 30320
rect 0 29656 800 29776
rect 0 29112 800 29232
rect 0 28568 800 28688
rect 67407 28568 68207 28688
rect 67407 28296 68207 28416
rect 0 28024 800 28144
rect 67407 28024 68207 28144
rect 67407 27752 68207 27872
rect 0 27480 800 27600
rect 67407 27480 68207 27600
rect 67407 27208 68207 27328
rect 0 26936 800 27056
rect 67407 26936 68207 27056
rect 67407 26664 68207 26784
rect 0 26392 800 26512
rect 67407 26392 68207 26512
rect 67407 26120 68207 26240
rect 0 25848 800 25968
rect 67407 25848 68207 25968
rect 67407 25576 68207 25696
rect 0 25304 800 25424
rect 67407 25304 68207 25424
rect 67407 25032 68207 25152
rect 0 24760 800 24880
rect 67407 24760 68207 24880
rect 67407 24488 68207 24608
rect 0 24216 800 24336
rect 67407 24216 68207 24336
rect 67407 23944 68207 24064
rect 0 23672 800 23792
rect 67407 23672 68207 23792
rect 67407 23400 68207 23520
rect 0 23128 800 23248
rect 67407 23128 68207 23248
rect 67407 22856 68207 22976
rect 0 22584 800 22704
rect 67407 22584 68207 22704
rect 67407 22312 68207 22432
rect 0 22040 800 22160
rect 67407 22040 68207 22160
rect 67407 21768 68207 21888
rect 0 21496 800 21616
rect 67407 21496 68207 21616
rect 67407 21224 68207 21344
rect 0 20952 800 21072
rect 67407 20952 68207 21072
rect 67407 20680 68207 20800
rect 0 20408 800 20528
rect 67407 20408 68207 20528
rect 67407 20136 68207 20256
rect 0 19864 800 19984
rect 67407 19864 68207 19984
rect 67407 19592 68207 19712
rect 0 19320 800 19440
rect 67407 19320 68207 19440
rect 67407 19048 68207 19168
rect 0 18776 800 18896
rect 67407 18776 68207 18896
rect 67407 18504 68207 18624
rect 0 18232 800 18352
rect 67407 18232 68207 18352
rect 67407 17960 68207 18080
rect 0 17688 800 17808
rect 67407 17688 68207 17808
rect 67407 17416 68207 17536
rect 0 17144 800 17264
rect 67407 17144 68207 17264
rect 67407 16872 68207 16992
rect 0 16600 800 16720
rect 67407 16600 68207 16720
rect 67407 16328 68207 16448
rect 0 16056 800 16176
rect 67407 16056 68207 16176
rect 67407 15784 68207 15904
rect 0 15512 800 15632
rect 67407 15512 68207 15632
rect 67407 15240 68207 15360
rect 0 14968 800 15088
rect 67407 14968 68207 15088
rect 67407 14696 68207 14816
rect 0 14424 800 14544
rect 67407 14424 68207 14544
rect 67407 14152 68207 14272
rect 0 13880 800 14000
rect 67407 13880 68207 14000
rect 67407 13608 68207 13728
rect 0 13336 800 13456
rect 67407 13336 68207 13456
rect 67407 13064 68207 13184
rect 0 12792 800 12912
rect 67407 12792 68207 12912
rect 67407 12520 68207 12640
rect 0 12248 800 12368
rect 67407 12248 68207 12368
rect 67407 11976 68207 12096
rect 0 11704 800 11824
rect 67407 11704 68207 11824
rect 67407 11432 68207 11552
rect 0 11160 800 11280
rect 67407 11160 68207 11280
rect 67407 10888 68207 11008
rect 0 10616 800 10736
rect 67407 10616 68207 10736
rect 67407 10344 68207 10464
rect 0 10072 800 10192
rect 67407 10072 68207 10192
rect 67407 9800 68207 9920
rect 0 9528 800 9648
rect 67407 9528 68207 9648
rect 67407 9256 68207 9376
rect 0 8984 800 9104
rect 67407 8984 68207 9104
rect 67407 8712 68207 8832
rect 0 8440 800 8560
rect 67407 8440 68207 8560
rect 0 7896 800 8016
rect 0 7352 800 7472
rect 0 6808 800 6928
rect 0 6264 800 6384
rect 0 5720 800 5840
rect 0 5176 800 5296
rect 0 4632 800 4752
rect 0 4088 800 4208
rect 0 3544 800 3664
rect 0 3000 800 3120
rect 0 2456 800 2576
rect 0 1912 800 2032
rect 0 1368 800 1488
rect 0 824 800 944
<< obsm3 >>
rect 800 35296 67407 35325
rect 880 35016 67407 35296
rect 800 34752 67407 35016
rect 880 34472 67407 34752
rect 800 34208 67407 34472
rect 880 33928 67407 34208
rect 800 33664 67407 33928
rect 880 33384 67407 33664
rect 800 33120 67407 33384
rect 880 32840 67407 33120
rect 800 32576 67407 32840
rect 880 32296 67407 32576
rect 800 32032 67407 32296
rect 880 31752 67407 32032
rect 800 31488 67407 31752
rect 880 31208 67407 31488
rect 800 30944 67407 31208
rect 880 30664 67407 30944
rect 800 30400 67407 30664
rect 880 30120 67407 30400
rect 800 29856 67407 30120
rect 880 29576 67407 29856
rect 800 29312 67407 29576
rect 880 29032 67407 29312
rect 800 28768 67407 29032
rect 880 28488 67327 28768
rect 800 28224 67327 28488
rect 880 27944 67327 28224
rect 800 27680 67327 27944
rect 880 27400 67327 27680
rect 800 27136 67327 27400
rect 880 26856 67327 27136
rect 800 26592 67327 26856
rect 880 26312 67327 26592
rect 800 26048 67327 26312
rect 880 25768 67327 26048
rect 800 25504 67327 25768
rect 880 25224 67327 25504
rect 800 24960 67327 25224
rect 880 24680 67327 24960
rect 800 24416 67327 24680
rect 880 24136 67327 24416
rect 800 23872 67327 24136
rect 880 23592 67327 23872
rect 800 23328 67327 23592
rect 880 23048 67327 23328
rect 800 22784 67327 23048
rect 880 22504 67327 22784
rect 800 22240 67327 22504
rect 880 21960 67327 22240
rect 800 21696 67327 21960
rect 880 21416 67327 21696
rect 800 21152 67327 21416
rect 880 20872 67327 21152
rect 800 20608 67327 20872
rect 880 20328 67327 20608
rect 800 20064 67327 20328
rect 880 19784 67327 20064
rect 800 19520 67327 19784
rect 880 19240 67327 19520
rect 800 18976 67327 19240
rect 880 18696 67327 18976
rect 800 18432 67327 18696
rect 880 18152 67327 18432
rect 800 17888 67327 18152
rect 880 17608 67327 17888
rect 800 17344 67327 17608
rect 880 17064 67327 17344
rect 800 16800 67327 17064
rect 880 16520 67327 16800
rect 800 16256 67327 16520
rect 880 15976 67327 16256
rect 800 15712 67327 15976
rect 880 15432 67327 15712
rect 800 15168 67327 15432
rect 880 14888 67327 15168
rect 800 14624 67327 14888
rect 880 14344 67327 14624
rect 800 14080 67327 14344
rect 880 13800 67327 14080
rect 800 13536 67327 13800
rect 880 13256 67327 13536
rect 800 12992 67327 13256
rect 880 12712 67327 12992
rect 800 12448 67327 12712
rect 880 12168 67327 12448
rect 800 11904 67327 12168
rect 880 11624 67327 11904
rect 800 11360 67327 11624
rect 880 11080 67327 11360
rect 800 10816 67327 11080
rect 880 10536 67327 10816
rect 800 10272 67327 10536
rect 880 9992 67327 10272
rect 800 9728 67327 9992
rect 880 9448 67327 9728
rect 800 9184 67327 9448
rect 880 8904 67327 9184
rect 800 8640 67327 8904
rect 880 8360 67327 8640
rect 800 8096 67407 8360
rect 880 7816 67407 8096
rect 800 7552 67407 7816
rect 880 7272 67407 7552
rect 800 7008 67407 7272
rect 880 6728 67407 7008
rect 800 6464 67407 6728
rect 880 6184 67407 6464
rect 800 5920 67407 6184
rect 880 5640 67407 5920
rect 800 5376 67407 5640
rect 880 5096 67407 5376
rect 800 4832 67407 5096
rect 880 4552 67407 4832
rect 800 4288 67407 4552
rect 880 4008 67407 4288
rect 800 3744 67407 4008
rect 880 3464 67407 3744
rect 800 3200 67407 3464
rect 880 2920 67407 3200
rect 800 2656 67407 2920
rect 880 2376 67407 2656
rect 800 2112 67407 2376
rect 880 1832 67407 2112
rect 800 1568 67407 1832
rect 880 1288 67407 1568
rect 800 1024 67407 1288
rect 880 744 67407 1024
rect 800 579 67407 744
<< metal4 >>
rect 9189 2128 9509 34864
rect 17434 2128 17754 34864
rect 25680 2128 26000 34864
rect 33925 2128 34245 34864
rect 42171 2128 42491 34864
rect 50416 2128 50736 34864
rect 58662 2128 58982 34864
rect 66907 2128 67227 34864
<< obsm4 >>
rect 2267 34944 66181 35325
rect 2267 2048 9109 34944
rect 9589 2048 17354 34944
rect 17834 2048 25600 34944
rect 26080 2048 33845 34944
rect 34325 2048 42091 34944
rect 42571 2048 50336 34944
rect 50816 2048 58582 34944
rect 59062 2048 66181 34944
rect 2267 715 66181 2048
<< obsm5 >>
rect 2876 4940 15156 12740
<< labels >>
rlabel metal3 s 67407 8984 68207 9104 6 becStatus[0]
port 1 nsew signal input
rlabel metal3 s 67407 9256 68207 9376 6 becStatus[1]
port 2 nsew signal input
rlabel metal3 s 67407 9528 68207 9648 6 becStatus[2]
port 3 nsew signal input
rlabel metal3 s 67407 9800 68207 9920 6 becStatus[3]
port 4 nsew signal input
rlabel metal2 s 4158 36551 4214 37351 6 data_in[0]
port 5 nsew signal input
rlabel metal2 s 22558 36551 22614 37351 6 data_in[100]
port 6 nsew signal input
rlabel metal2 s 22742 36551 22798 37351 6 data_in[101]
port 7 nsew signal input
rlabel metal2 s 22926 36551 22982 37351 6 data_in[102]
port 8 nsew signal input
rlabel metal2 s 23110 36551 23166 37351 6 data_in[103]
port 9 nsew signal input
rlabel metal2 s 23294 36551 23350 37351 6 data_in[104]
port 10 nsew signal input
rlabel metal2 s 23478 36551 23534 37351 6 data_in[105]
port 11 nsew signal input
rlabel metal2 s 23662 36551 23718 37351 6 data_in[106]
port 12 nsew signal input
rlabel metal2 s 23846 36551 23902 37351 6 data_in[107]
port 13 nsew signal input
rlabel metal2 s 24030 36551 24086 37351 6 data_in[108]
port 14 nsew signal input
rlabel metal2 s 24214 36551 24270 37351 6 data_in[109]
port 15 nsew signal input
rlabel metal2 s 5998 36551 6054 37351 6 data_in[10]
port 16 nsew signal input
rlabel metal2 s 24398 36551 24454 37351 6 data_in[110]
port 17 nsew signal input
rlabel metal2 s 24582 36551 24638 37351 6 data_in[111]
port 18 nsew signal input
rlabel metal2 s 24766 36551 24822 37351 6 data_in[112]
port 19 nsew signal input
rlabel metal2 s 24950 36551 25006 37351 6 data_in[113]
port 20 nsew signal input
rlabel metal2 s 25134 36551 25190 37351 6 data_in[114]
port 21 nsew signal input
rlabel metal2 s 25318 36551 25374 37351 6 data_in[115]
port 22 nsew signal input
rlabel metal2 s 25502 36551 25558 37351 6 data_in[116]
port 23 nsew signal input
rlabel metal2 s 25686 36551 25742 37351 6 data_in[117]
port 24 nsew signal input
rlabel metal2 s 25870 36551 25926 37351 6 data_in[118]
port 25 nsew signal input
rlabel metal2 s 26054 36551 26110 37351 6 data_in[119]
port 26 nsew signal input
rlabel metal2 s 6182 36551 6238 37351 6 data_in[11]
port 27 nsew signal input
rlabel metal2 s 26238 36551 26294 37351 6 data_in[120]
port 28 nsew signal input
rlabel metal2 s 26422 36551 26478 37351 6 data_in[121]
port 29 nsew signal input
rlabel metal2 s 26606 36551 26662 37351 6 data_in[122]
port 30 nsew signal input
rlabel metal2 s 26790 36551 26846 37351 6 data_in[123]
port 31 nsew signal input
rlabel metal2 s 26974 36551 27030 37351 6 data_in[124]
port 32 nsew signal input
rlabel metal2 s 27158 36551 27214 37351 6 data_in[125]
port 33 nsew signal input
rlabel metal2 s 27342 36551 27398 37351 6 data_in[126]
port 34 nsew signal input
rlabel metal2 s 27526 36551 27582 37351 6 data_in[127]
port 35 nsew signal input
rlabel metal2 s 27710 36551 27766 37351 6 data_in[128]
port 36 nsew signal input
rlabel metal2 s 27894 36551 27950 37351 6 data_in[129]
port 37 nsew signal input
rlabel metal2 s 6366 36551 6422 37351 6 data_in[12]
port 38 nsew signal input
rlabel metal2 s 28078 36551 28134 37351 6 data_in[130]
port 39 nsew signal input
rlabel metal2 s 28262 36551 28318 37351 6 data_in[131]
port 40 nsew signal input
rlabel metal2 s 28446 36551 28502 37351 6 data_in[132]
port 41 nsew signal input
rlabel metal2 s 28630 36551 28686 37351 6 data_in[133]
port 42 nsew signal input
rlabel metal2 s 28814 36551 28870 37351 6 data_in[134]
port 43 nsew signal input
rlabel metal2 s 28998 36551 29054 37351 6 data_in[135]
port 44 nsew signal input
rlabel metal2 s 29182 36551 29238 37351 6 data_in[136]
port 45 nsew signal input
rlabel metal2 s 29366 36551 29422 37351 6 data_in[137]
port 46 nsew signal input
rlabel metal2 s 29550 36551 29606 37351 6 data_in[138]
port 47 nsew signal input
rlabel metal2 s 29734 36551 29790 37351 6 data_in[139]
port 48 nsew signal input
rlabel metal2 s 6550 36551 6606 37351 6 data_in[13]
port 49 nsew signal input
rlabel metal2 s 29918 36551 29974 37351 6 data_in[140]
port 50 nsew signal input
rlabel metal2 s 30102 36551 30158 37351 6 data_in[141]
port 51 nsew signal input
rlabel metal2 s 30286 36551 30342 37351 6 data_in[142]
port 52 nsew signal input
rlabel metal2 s 30470 36551 30526 37351 6 data_in[143]
port 53 nsew signal input
rlabel metal2 s 30654 36551 30710 37351 6 data_in[144]
port 54 nsew signal input
rlabel metal2 s 30838 36551 30894 37351 6 data_in[145]
port 55 nsew signal input
rlabel metal2 s 31022 36551 31078 37351 6 data_in[146]
port 56 nsew signal input
rlabel metal2 s 31206 36551 31262 37351 6 data_in[147]
port 57 nsew signal input
rlabel metal2 s 31390 36551 31446 37351 6 data_in[148]
port 58 nsew signal input
rlabel metal2 s 31574 36551 31630 37351 6 data_in[149]
port 59 nsew signal input
rlabel metal2 s 6734 36551 6790 37351 6 data_in[14]
port 60 nsew signal input
rlabel metal2 s 31758 36551 31814 37351 6 data_in[150]
port 61 nsew signal input
rlabel metal2 s 31942 36551 31998 37351 6 data_in[151]
port 62 nsew signal input
rlabel metal2 s 32126 36551 32182 37351 6 data_in[152]
port 63 nsew signal input
rlabel metal2 s 32310 36551 32366 37351 6 data_in[153]
port 64 nsew signal input
rlabel metal2 s 32494 36551 32550 37351 6 data_in[154]
port 65 nsew signal input
rlabel metal2 s 32678 36551 32734 37351 6 data_in[155]
port 66 nsew signal input
rlabel metal2 s 32862 36551 32918 37351 6 data_in[156]
port 67 nsew signal input
rlabel metal2 s 33046 36551 33102 37351 6 data_in[157]
port 68 nsew signal input
rlabel metal2 s 33230 36551 33286 37351 6 data_in[158]
port 69 nsew signal input
rlabel metal2 s 33414 36551 33470 37351 6 data_in[159]
port 70 nsew signal input
rlabel metal2 s 6918 36551 6974 37351 6 data_in[15]
port 71 nsew signal input
rlabel metal2 s 33598 36551 33654 37351 6 data_in[160]
port 72 nsew signal input
rlabel metal2 s 33782 36551 33838 37351 6 data_in[161]
port 73 nsew signal input
rlabel metal2 s 33966 36551 34022 37351 6 data_in[162]
port 74 nsew signal input
rlabel metal2 s 7102 36551 7158 37351 6 data_in[16]
port 75 nsew signal input
rlabel metal2 s 7286 36551 7342 37351 6 data_in[17]
port 76 nsew signal input
rlabel metal2 s 7470 36551 7526 37351 6 data_in[18]
port 77 nsew signal input
rlabel metal2 s 7654 36551 7710 37351 6 data_in[19]
port 78 nsew signal input
rlabel metal2 s 4342 36551 4398 37351 6 data_in[1]
port 79 nsew signal input
rlabel metal2 s 7838 36551 7894 37351 6 data_in[20]
port 80 nsew signal input
rlabel metal2 s 8022 36551 8078 37351 6 data_in[21]
port 81 nsew signal input
rlabel metal2 s 8206 36551 8262 37351 6 data_in[22]
port 82 nsew signal input
rlabel metal2 s 8390 36551 8446 37351 6 data_in[23]
port 83 nsew signal input
rlabel metal2 s 8574 36551 8630 37351 6 data_in[24]
port 84 nsew signal input
rlabel metal2 s 8758 36551 8814 37351 6 data_in[25]
port 85 nsew signal input
rlabel metal2 s 8942 36551 8998 37351 6 data_in[26]
port 86 nsew signal input
rlabel metal2 s 9126 36551 9182 37351 6 data_in[27]
port 87 nsew signal input
rlabel metal2 s 9310 36551 9366 37351 6 data_in[28]
port 88 nsew signal input
rlabel metal2 s 9494 36551 9550 37351 6 data_in[29]
port 89 nsew signal input
rlabel metal2 s 4526 36551 4582 37351 6 data_in[2]
port 90 nsew signal input
rlabel metal2 s 9678 36551 9734 37351 6 data_in[30]
port 91 nsew signal input
rlabel metal2 s 9862 36551 9918 37351 6 data_in[31]
port 92 nsew signal input
rlabel metal2 s 10046 36551 10102 37351 6 data_in[32]
port 93 nsew signal input
rlabel metal2 s 10230 36551 10286 37351 6 data_in[33]
port 94 nsew signal input
rlabel metal2 s 10414 36551 10470 37351 6 data_in[34]
port 95 nsew signal input
rlabel metal2 s 10598 36551 10654 37351 6 data_in[35]
port 96 nsew signal input
rlabel metal2 s 10782 36551 10838 37351 6 data_in[36]
port 97 nsew signal input
rlabel metal2 s 10966 36551 11022 37351 6 data_in[37]
port 98 nsew signal input
rlabel metal2 s 11150 36551 11206 37351 6 data_in[38]
port 99 nsew signal input
rlabel metal2 s 11334 36551 11390 37351 6 data_in[39]
port 100 nsew signal input
rlabel metal2 s 4710 36551 4766 37351 6 data_in[3]
port 101 nsew signal input
rlabel metal2 s 11518 36551 11574 37351 6 data_in[40]
port 102 nsew signal input
rlabel metal2 s 11702 36551 11758 37351 6 data_in[41]
port 103 nsew signal input
rlabel metal2 s 11886 36551 11942 37351 6 data_in[42]
port 104 nsew signal input
rlabel metal2 s 12070 36551 12126 37351 6 data_in[43]
port 105 nsew signal input
rlabel metal2 s 12254 36551 12310 37351 6 data_in[44]
port 106 nsew signal input
rlabel metal2 s 12438 36551 12494 37351 6 data_in[45]
port 107 nsew signal input
rlabel metal2 s 12622 36551 12678 37351 6 data_in[46]
port 108 nsew signal input
rlabel metal2 s 12806 36551 12862 37351 6 data_in[47]
port 109 nsew signal input
rlabel metal2 s 12990 36551 13046 37351 6 data_in[48]
port 110 nsew signal input
rlabel metal2 s 13174 36551 13230 37351 6 data_in[49]
port 111 nsew signal input
rlabel metal2 s 4894 36551 4950 37351 6 data_in[4]
port 112 nsew signal input
rlabel metal2 s 13358 36551 13414 37351 6 data_in[50]
port 113 nsew signal input
rlabel metal2 s 13542 36551 13598 37351 6 data_in[51]
port 114 nsew signal input
rlabel metal2 s 13726 36551 13782 37351 6 data_in[52]
port 115 nsew signal input
rlabel metal2 s 13910 36551 13966 37351 6 data_in[53]
port 116 nsew signal input
rlabel metal2 s 14094 36551 14150 37351 6 data_in[54]
port 117 nsew signal input
rlabel metal2 s 14278 36551 14334 37351 6 data_in[55]
port 118 nsew signal input
rlabel metal2 s 14462 36551 14518 37351 6 data_in[56]
port 119 nsew signal input
rlabel metal2 s 14646 36551 14702 37351 6 data_in[57]
port 120 nsew signal input
rlabel metal2 s 14830 36551 14886 37351 6 data_in[58]
port 121 nsew signal input
rlabel metal2 s 15014 36551 15070 37351 6 data_in[59]
port 122 nsew signal input
rlabel metal2 s 5078 36551 5134 37351 6 data_in[5]
port 123 nsew signal input
rlabel metal2 s 15198 36551 15254 37351 6 data_in[60]
port 124 nsew signal input
rlabel metal2 s 15382 36551 15438 37351 6 data_in[61]
port 125 nsew signal input
rlabel metal2 s 15566 36551 15622 37351 6 data_in[62]
port 126 nsew signal input
rlabel metal2 s 15750 36551 15806 37351 6 data_in[63]
port 127 nsew signal input
rlabel metal2 s 15934 36551 15990 37351 6 data_in[64]
port 128 nsew signal input
rlabel metal2 s 16118 36551 16174 37351 6 data_in[65]
port 129 nsew signal input
rlabel metal2 s 16302 36551 16358 37351 6 data_in[66]
port 130 nsew signal input
rlabel metal2 s 16486 36551 16542 37351 6 data_in[67]
port 131 nsew signal input
rlabel metal2 s 16670 36551 16726 37351 6 data_in[68]
port 132 nsew signal input
rlabel metal2 s 16854 36551 16910 37351 6 data_in[69]
port 133 nsew signal input
rlabel metal2 s 5262 36551 5318 37351 6 data_in[6]
port 134 nsew signal input
rlabel metal2 s 17038 36551 17094 37351 6 data_in[70]
port 135 nsew signal input
rlabel metal2 s 17222 36551 17278 37351 6 data_in[71]
port 136 nsew signal input
rlabel metal2 s 17406 36551 17462 37351 6 data_in[72]
port 137 nsew signal input
rlabel metal2 s 17590 36551 17646 37351 6 data_in[73]
port 138 nsew signal input
rlabel metal2 s 17774 36551 17830 37351 6 data_in[74]
port 139 nsew signal input
rlabel metal2 s 17958 36551 18014 37351 6 data_in[75]
port 140 nsew signal input
rlabel metal2 s 18142 36551 18198 37351 6 data_in[76]
port 141 nsew signal input
rlabel metal2 s 18326 36551 18382 37351 6 data_in[77]
port 142 nsew signal input
rlabel metal2 s 18510 36551 18566 37351 6 data_in[78]
port 143 nsew signal input
rlabel metal2 s 18694 36551 18750 37351 6 data_in[79]
port 144 nsew signal input
rlabel metal2 s 5446 36551 5502 37351 6 data_in[7]
port 145 nsew signal input
rlabel metal2 s 18878 36551 18934 37351 6 data_in[80]
port 146 nsew signal input
rlabel metal2 s 19062 36551 19118 37351 6 data_in[81]
port 147 nsew signal input
rlabel metal2 s 19246 36551 19302 37351 6 data_in[82]
port 148 nsew signal input
rlabel metal2 s 19430 36551 19486 37351 6 data_in[83]
port 149 nsew signal input
rlabel metal2 s 19614 36551 19670 37351 6 data_in[84]
port 150 nsew signal input
rlabel metal2 s 19798 36551 19854 37351 6 data_in[85]
port 151 nsew signal input
rlabel metal2 s 19982 36551 20038 37351 6 data_in[86]
port 152 nsew signal input
rlabel metal2 s 20166 36551 20222 37351 6 data_in[87]
port 153 nsew signal input
rlabel metal2 s 20350 36551 20406 37351 6 data_in[88]
port 154 nsew signal input
rlabel metal2 s 20534 36551 20590 37351 6 data_in[89]
port 155 nsew signal input
rlabel metal2 s 5630 36551 5686 37351 6 data_in[8]
port 156 nsew signal input
rlabel metal2 s 20718 36551 20774 37351 6 data_in[90]
port 157 nsew signal input
rlabel metal2 s 20902 36551 20958 37351 6 data_in[91]
port 158 nsew signal input
rlabel metal2 s 21086 36551 21142 37351 6 data_in[92]
port 159 nsew signal input
rlabel metal2 s 21270 36551 21326 37351 6 data_in[93]
port 160 nsew signal input
rlabel metal2 s 21454 36551 21510 37351 6 data_in[94]
port 161 nsew signal input
rlabel metal2 s 21638 36551 21694 37351 6 data_in[95]
port 162 nsew signal input
rlabel metal2 s 21822 36551 21878 37351 6 data_in[96]
port 163 nsew signal input
rlabel metal2 s 22006 36551 22062 37351 6 data_in[97]
port 164 nsew signal input
rlabel metal2 s 22190 36551 22246 37351 6 data_in[98]
port 165 nsew signal input
rlabel metal2 s 22374 36551 22430 37351 6 data_in[99]
port 166 nsew signal input
rlabel metal2 s 5814 36551 5870 37351 6 data_in[9]
port 167 nsew signal input
rlabel metal2 s 34150 36551 34206 37351 6 data_out[0]
port 168 nsew signal output
rlabel metal2 s 52550 36551 52606 37351 6 data_out[100]
port 169 nsew signal output
rlabel metal2 s 52734 36551 52790 37351 6 data_out[101]
port 170 nsew signal output
rlabel metal2 s 52918 36551 52974 37351 6 data_out[102]
port 171 nsew signal output
rlabel metal2 s 53102 36551 53158 37351 6 data_out[103]
port 172 nsew signal output
rlabel metal2 s 53286 36551 53342 37351 6 data_out[104]
port 173 nsew signal output
rlabel metal2 s 53470 36551 53526 37351 6 data_out[105]
port 174 nsew signal output
rlabel metal2 s 53654 36551 53710 37351 6 data_out[106]
port 175 nsew signal output
rlabel metal2 s 53838 36551 53894 37351 6 data_out[107]
port 176 nsew signal output
rlabel metal2 s 54022 36551 54078 37351 6 data_out[108]
port 177 nsew signal output
rlabel metal2 s 54206 36551 54262 37351 6 data_out[109]
port 178 nsew signal output
rlabel metal2 s 35990 36551 36046 37351 6 data_out[10]
port 179 nsew signal output
rlabel metal2 s 54390 36551 54446 37351 6 data_out[110]
port 180 nsew signal output
rlabel metal2 s 54574 36551 54630 37351 6 data_out[111]
port 181 nsew signal output
rlabel metal2 s 54758 36551 54814 37351 6 data_out[112]
port 182 nsew signal output
rlabel metal2 s 54942 36551 54998 37351 6 data_out[113]
port 183 nsew signal output
rlabel metal2 s 55126 36551 55182 37351 6 data_out[114]
port 184 nsew signal output
rlabel metal2 s 55310 36551 55366 37351 6 data_out[115]
port 185 nsew signal output
rlabel metal2 s 55494 36551 55550 37351 6 data_out[116]
port 186 nsew signal output
rlabel metal2 s 55678 36551 55734 37351 6 data_out[117]
port 187 nsew signal output
rlabel metal2 s 55862 36551 55918 37351 6 data_out[118]
port 188 nsew signal output
rlabel metal2 s 56046 36551 56102 37351 6 data_out[119]
port 189 nsew signal output
rlabel metal2 s 36174 36551 36230 37351 6 data_out[11]
port 190 nsew signal output
rlabel metal2 s 56230 36551 56286 37351 6 data_out[120]
port 191 nsew signal output
rlabel metal2 s 56414 36551 56470 37351 6 data_out[121]
port 192 nsew signal output
rlabel metal2 s 56598 36551 56654 37351 6 data_out[122]
port 193 nsew signal output
rlabel metal2 s 56782 36551 56838 37351 6 data_out[123]
port 194 nsew signal output
rlabel metal2 s 56966 36551 57022 37351 6 data_out[124]
port 195 nsew signal output
rlabel metal2 s 57150 36551 57206 37351 6 data_out[125]
port 196 nsew signal output
rlabel metal2 s 57334 36551 57390 37351 6 data_out[126]
port 197 nsew signal output
rlabel metal2 s 57518 36551 57574 37351 6 data_out[127]
port 198 nsew signal output
rlabel metal2 s 57702 36551 57758 37351 6 data_out[128]
port 199 nsew signal output
rlabel metal2 s 57886 36551 57942 37351 6 data_out[129]
port 200 nsew signal output
rlabel metal2 s 36358 36551 36414 37351 6 data_out[12]
port 201 nsew signal output
rlabel metal2 s 58070 36551 58126 37351 6 data_out[130]
port 202 nsew signal output
rlabel metal2 s 58254 36551 58310 37351 6 data_out[131]
port 203 nsew signal output
rlabel metal2 s 58438 36551 58494 37351 6 data_out[132]
port 204 nsew signal output
rlabel metal2 s 58622 36551 58678 37351 6 data_out[133]
port 205 nsew signal output
rlabel metal2 s 58806 36551 58862 37351 6 data_out[134]
port 206 nsew signal output
rlabel metal2 s 58990 36551 59046 37351 6 data_out[135]
port 207 nsew signal output
rlabel metal2 s 59174 36551 59230 37351 6 data_out[136]
port 208 nsew signal output
rlabel metal2 s 59358 36551 59414 37351 6 data_out[137]
port 209 nsew signal output
rlabel metal2 s 59542 36551 59598 37351 6 data_out[138]
port 210 nsew signal output
rlabel metal2 s 59726 36551 59782 37351 6 data_out[139]
port 211 nsew signal output
rlabel metal2 s 36542 36551 36598 37351 6 data_out[13]
port 212 nsew signal output
rlabel metal2 s 59910 36551 59966 37351 6 data_out[140]
port 213 nsew signal output
rlabel metal2 s 60094 36551 60150 37351 6 data_out[141]
port 214 nsew signal output
rlabel metal2 s 60278 36551 60334 37351 6 data_out[142]
port 215 nsew signal output
rlabel metal2 s 60462 36551 60518 37351 6 data_out[143]
port 216 nsew signal output
rlabel metal2 s 60646 36551 60702 37351 6 data_out[144]
port 217 nsew signal output
rlabel metal2 s 60830 36551 60886 37351 6 data_out[145]
port 218 nsew signal output
rlabel metal2 s 61014 36551 61070 37351 6 data_out[146]
port 219 nsew signal output
rlabel metal2 s 61198 36551 61254 37351 6 data_out[147]
port 220 nsew signal output
rlabel metal2 s 61382 36551 61438 37351 6 data_out[148]
port 221 nsew signal output
rlabel metal2 s 61566 36551 61622 37351 6 data_out[149]
port 222 nsew signal output
rlabel metal2 s 36726 36551 36782 37351 6 data_out[14]
port 223 nsew signal output
rlabel metal2 s 61750 36551 61806 37351 6 data_out[150]
port 224 nsew signal output
rlabel metal2 s 61934 36551 61990 37351 6 data_out[151]
port 225 nsew signal output
rlabel metal2 s 62118 36551 62174 37351 6 data_out[152]
port 226 nsew signal output
rlabel metal2 s 62302 36551 62358 37351 6 data_out[153]
port 227 nsew signal output
rlabel metal2 s 62486 36551 62542 37351 6 data_out[154]
port 228 nsew signal output
rlabel metal2 s 62670 36551 62726 37351 6 data_out[155]
port 229 nsew signal output
rlabel metal2 s 62854 36551 62910 37351 6 data_out[156]
port 230 nsew signal output
rlabel metal2 s 63038 36551 63094 37351 6 data_out[157]
port 231 nsew signal output
rlabel metal2 s 63222 36551 63278 37351 6 data_out[158]
port 232 nsew signal output
rlabel metal2 s 63406 36551 63462 37351 6 data_out[159]
port 233 nsew signal output
rlabel metal2 s 36910 36551 36966 37351 6 data_out[15]
port 234 nsew signal output
rlabel metal2 s 63590 36551 63646 37351 6 data_out[160]
port 235 nsew signal output
rlabel metal2 s 63774 36551 63830 37351 6 data_out[161]
port 236 nsew signal output
rlabel metal2 s 63958 36551 64014 37351 6 data_out[162]
port 237 nsew signal output
rlabel metal2 s 37094 36551 37150 37351 6 data_out[16]
port 238 nsew signal output
rlabel metal2 s 37278 36551 37334 37351 6 data_out[17]
port 239 nsew signal output
rlabel metal2 s 37462 36551 37518 37351 6 data_out[18]
port 240 nsew signal output
rlabel metal2 s 37646 36551 37702 37351 6 data_out[19]
port 241 nsew signal output
rlabel metal2 s 34334 36551 34390 37351 6 data_out[1]
port 242 nsew signal output
rlabel metal2 s 37830 36551 37886 37351 6 data_out[20]
port 243 nsew signal output
rlabel metal2 s 38014 36551 38070 37351 6 data_out[21]
port 244 nsew signal output
rlabel metal2 s 38198 36551 38254 37351 6 data_out[22]
port 245 nsew signal output
rlabel metal2 s 38382 36551 38438 37351 6 data_out[23]
port 246 nsew signal output
rlabel metal2 s 38566 36551 38622 37351 6 data_out[24]
port 247 nsew signal output
rlabel metal2 s 38750 36551 38806 37351 6 data_out[25]
port 248 nsew signal output
rlabel metal2 s 38934 36551 38990 37351 6 data_out[26]
port 249 nsew signal output
rlabel metal2 s 39118 36551 39174 37351 6 data_out[27]
port 250 nsew signal output
rlabel metal2 s 39302 36551 39358 37351 6 data_out[28]
port 251 nsew signal output
rlabel metal2 s 39486 36551 39542 37351 6 data_out[29]
port 252 nsew signal output
rlabel metal2 s 34518 36551 34574 37351 6 data_out[2]
port 253 nsew signal output
rlabel metal2 s 39670 36551 39726 37351 6 data_out[30]
port 254 nsew signal output
rlabel metal2 s 39854 36551 39910 37351 6 data_out[31]
port 255 nsew signal output
rlabel metal2 s 40038 36551 40094 37351 6 data_out[32]
port 256 nsew signal output
rlabel metal2 s 40222 36551 40278 37351 6 data_out[33]
port 257 nsew signal output
rlabel metal2 s 40406 36551 40462 37351 6 data_out[34]
port 258 nsew signal output
rlabel metal2 s 40590 36551 40646 37351 6 data_out[35]
port 259 nsew signal output
rlabel metal2 s 40774 36551 40830 37351 6 data_out[36]
port 260 nsew signal output
rlabel metal2 s 40958 36551 41014 37351 6 data_out[37]
port 261 nsew signal output
rlabel metal2 s 41142 36551 41198 37351 6 data_out[38]
port 262 nsew signal output
rlabel metal2 s 41326 36551 41382 37351 6 data_out[39]
port 263 nsew signal output
rlabel metal2 s 34702 36551 34758 37351 6 data_out[3]
port 264 nsew signal output
rlabel metal2 s 41510 36551 41566 37351 6 data_out[40]
port 265 nsew signal output
rlabel metal2 s 41694 36551 41750 37351 6 data_out[41]
port 266 nsew signal output
rlabel metal2 s 41878 36551 41934 37351 6 data_out[42]
port 267 nsew signal output
rlabel metal2 s 42062 36551 42118 37351 6 data_out[43]
port 268 nsew signal output
rlabel metal2 s 42246 36551 42302 37351 6 data_out[44]
port 269 nsew signal output
rlabel metal2 s 42430 36551 42486 37351 6 data_out[45]
port 270 nsew signal output
rlabel metal2 s 42614 36551 42670 37351 6 data_out[46]
port 271 nsew signal output
rlabel metal2 s 42798 36551 42854 37351 6 data_out[47]
port 272 nsew signal output
rlabel metal2 s 42982 36551 43038 37351 6 data_out[48]
port 273 nsew signal output
rlabel metal2 s 43166 36551 43222 37351 6 data_out[49]
port 274 nsew signal output
rlabel metal2 s 34886 36551 34942 37351 6 data_out[4]
port 275 nsew signal output
rlabel metal2 s 43350 36551 43406 37351 6 data_out[50]
port 276 nsew signal output
rlabel metal2 s 43534 36551 43590 37351 6 data_out[51]
port 277 nsew signal output
rlabel metal2 s 43718 36551 43774 37351 6 data_out[52]
port 278 nsew signal output
rlabel metal2 s 43902 36551 43958 37351 6 data_out[53]
port 279 nsew signal output
rlabel metal2 s 44086 36551 44142 37351 6 data_out[54]
port 280 nsew signal output
rlabel metal2 s 44270 36551 44326 37351 6 data_out[55]
port 281 nsew signal output
rlabel metal2 s 44454 36551 44510 37351 6 data_out[56]
port 282 nsew signal output
rlabel metal2 s 44638 36551 44694 37351 6 data_out[57]
port 283 nsew signal output
rlabel metal2 s 44822 36551 44878 37351 6 data_out[58]
port 284 nsew signal output
rlabel metal2 s 45006 36551 45062 37351 6 data_out[59]
port 285 nsew signal output
rlabel metal2 s 35070 36551 35126 37351 6 data_out[5]
port 286 nsew signal output
rlabel metal2 s 45190 36551 45246 37351 6 data_out[60]
port 287 nsew signal output
rlabel metal2 s 45374 36551 45430 37351 6 data_out[61]
port 288 nsew signal output
rlabel metal2 s 45558 36551 45614 37351 6 data_out[62]
port 289 nsew signal output
rlabel metal2 s 45742 36551 45798 37351 6 data_out[63]
port 290 nsew signal output
rlabel metal2 s 45926 36551 45982 37351 6 data_out[64]
port 291 nsew signal output
rlabel metal2 s 46110 36551 46166 37351 6 data_out[65]
port 292 nsew signal output
rlabel metal2 s 46294 36551 46350 37351 6 data_out[66]
port 293 nsew signal output
rlabel metal2 s 46478 36551 46534 37351 6 data_out[67]
port 294 nsew signal output
rlabel metal2 s 46662 36551 46718 37351 6 data_out[68]
port 295 nsew signal output
rlabel metal2 s 46846 36551 46902 37351 6 data_out[69]
port 296 nsew signal output
rlabel metal2 s 35254 36551 35310 37351 6 data_out[6]
port 297 nsew signal output
rlabel metal2 s 47030 36551 47086 37351 6 data_out[70]
port 298 nsew signal output
rlabel metal2 s 47214 36551 47270 37351 6 data_out[71]
port 299 nsew signal output
rlabel metal2 s 47398 36551 47454 37351 6 data_out[72]
port 300 nsew signal output
rlabel metal2 s 47582 36551 47638 37351 6 data_out[73]
port 301 nsew signal output
rlabel metal2 s 47766 36551 47822 37351 6 data_out[74]
port 302 nsew signal output
rlabel metal2 s 47950 36551 48006 37351 6 data_out[75]
port 303 nsew signal output
rlabel metal2 s 48134 36551 48190 37351 6 data_out[76]
port 304 nsew signal output
rlabel metal2 s 48318 36551 48374 37351 6 data_out[77]
port 305 nsew signal output
rlabel metal2 s 48502 36551 48558 37351 6 data_out[78]
port 306 nsew signal output
rlabel metal2 s 48686 36551 48742 37351 6 data_out[79]
port 307 nsew signal output
rlabel metal2 s 35438 36551 35494 37351 6 data_out[7]
port 308 nsew signal output
rlabel metal2 s 48870 36551 48926 37351 6 data_out[80]
port 309 nsew signal output
rlabel metal2 s 49054 36551 49110 37351 6 data_out[81]
port 310 nsew signal output
rlabel metal2 s 49238 36551 49294 37351 6 data_out[82]
port 311 nsew signal output
rlabel metal2 s 49422 36551 49478 37351 6 data_out[83]
port 312 nsew signal output
rlabel metal2 s 49606 36551 49662 37351 6 data_out[84]
port 313 nsew signal output
rlabel metal2 s 49790 36551 49846 37351 6 data_out[85]
port 314 nsew signal output
rlabel metal2 s 49974 36551 50030 37351 6 data_out[86]
port 315 nsew signal output
rlabel metal2 s 50158 36551 50214 37351 6 data_out[87]
port 316 nsew signal output
rlabel metal2 s 50342 36551 50398 37351 6 data_out[88]
port 317 nsew signal output
rlabel metal2 s 50526 36551 50582 37351 6 data_out[89]
port 318 nsew signal output
rlabel metal2 s 35622 36551 35678 37351 6 data_out[8]
port 319 nsew signal output
rlabel metal2 s 50710 36551 50766 37351 6 data_out[90]
port 320 nsew signal output
rlabel metal2 s 50894 36551 50950 37351 6 data_out[91]
port 321 nsew signal output
rlabel metal2 s 51078 36551 51134 37351 6 data_out[92]
port 322 nsew signal output
rlabel metal2 s 51262 36551 51318 37351 6 data_out[93]
port 323 nsew signal output
rlabel metal2 s 51446 36551 51502 37351 6 data_out[94]
port 324 nsew signal output
rlabel metal2 s 51630 36551 51686 37351 6 data_out[95]
port 325 nsew signal output
rlabel metal2 s 51814 36551 51870 37351 6 data_out[96]
port 326 nsew signal output
rlabel metal2 s 51998 36551 52054 37351 6 data_out[97]
port 327 nsew signal output
rlabel metal2 s 52182 36551 52238 37351 6 data_out[98]
port 328 nsew signal output
rlabel metal2 s 52366 36551 52422 37351 6 data_out[99]
port 329 nsew signal output
rlabel metal2 s 35806 36551 35862 37351 6 data_out[9]
port 330 nsew signal output
rlabel metal3 s 0 2456 800 2576 6 ki
port 331 nsew signal output
rlabel metal2 s 10782 0 10838 800 6 la_data_in[0]
port 332 nsew signal input
rlabel metal2 s 29182 0 29238 800 6 la_data_in[100]
port 333 nsew signal input
rlabel metal2 s 29366 0 29422 800 6 la_data_in[101]
port 334 nsew signal input
rlabel metal2 s 29550 0 29606 800 6 la_data_in[102]
port 335 nsew signal input
rlabel metal2 s 29734 0 29790 800 6 la_data_in[103]
port 336 nsew signal input
rlabel metal2 s 29918 0 29974 800 6 la_data_in[104]
port 337 nsew signal input
rlabel metal2 s 30102 0 30158 800 6 la_data_in[105]
port 338 nsew signal input
rlabel metal2 s 30286 0 30342 800 6 la_data_in[106]
port 339 nsew signal input
rlabel metal2 s 30470 0 30526 800 6 la_data_in[107]
port 340 nsew signal input
rlabel metal2 s 30654 0 30710 800 6 la_data_in[108]
port 341 nsew signal input
rlabel metal2 s 30838 0 30894 800 6 la_data_in[109]
port 342 nsew signal input
rlabel metal2 s 12622 0 12678 800 6 la_data_in[10]
port 343 nsew signal input
rlabel metal2 s 31022 0 31078 800 6 la_data_in[110]
port 344 nsew signal input
rlabel metal2 s 31206 0 31262 800 6 la_data_in[111]
port 345 nsew signal input
rlabel metal2 s 31390 0 31446 800 6 la_data_in[112]
port 346 nsew signal input
rlabel metal2 s 31574 0 31630 800 6 la_data_in[113]
port 347 nsew signal input
rlabel metal2 s 31758 0 31814 800 6 la_data_in[114]
port 348 nsew signal input
rlabel metal2 s 31942 0 31998 800 6 la_data_in[115]
port 349 nsew signal input
rlabel metal2 s 32126 0 32182 800 6 la_data_in[116]
port 350 nsew signal input
rlabel metal2 s 32310 0 32366 800 6 la_data_in[117]
port 351 nsew signal input
rlabel metal2 s 32494 0 32550 800 6 la_data_in[118]
port 352 nsew signal input
rlabel metal2 s 32678 0 32734 800 6 la_data_in[119]
port 353 nsew signal input
rlabel metal2 s 12806 0 12862 800 6 la_data_in[11]
port 354 nsew signal input
rlabel metal2 s 32862 0 32918 800 6 la_data_in[120]
port 355 nsew signal input
rlabel metal2 s 33046 0 33102 800 6 la_data_in[121]
port 356 nsew signal input
rlabel metal2 s 33230 0 33286 800 6 la_data_in[122]
port 357 nsew signal input
rlabel metal2 s 33414 0 33470 800 6 la_data_in[123]
port 358 nsew signal input
rlabel metal2 s 33598 0 33654 800 6 la_data_in[124]
port 359 nsew signal input
rlabel metal2 s 33782 0 33838 800 6 la_data_in[125]
port 360 nsew signal input
rlabel metal2 s 33966 0 34022 800 6 la_data_in[126]
port 361 nsew signal input
rlabel metal2 s 34150 0 34206 800 6 la_data_in[127]
port 362 nsew signal input
rlabel metal2 s 12990 0 13046 800 6 la_data_in[12]
port 363 nsew signal input
rlabel metal2 s 13174 0 13230 800 6 la_data_in[13]
port 364 nsew signal input
rlabel metal2 s 13358 0 13414 800 6 la_data_in[14]
port 365 nsew signal input
rlabel metal2 s 13542 0 13598 800 6 la_data_in[15]
port 366 nsew signal input
rlabel metal2 s 13726 0 13782 800 6 la_data_in[16]
port 367 nsew signal input
rlabel metal2 s 13910 0 13966 800 6 la_data_in[17]
port 368 nsew signal input
rlabel metal2 s 14094 0 14150 800 6 la_data_in[18]
port 369 nsew signal input
rlabel metal2 s 14278 0 14334 800 6 la_data_in[19]
port 370 nsew signal input
rlabel metal2 s 10966 0 11022 800 6 la_data_in[1]
port 371 nsew signal input
rlabel metal2 s 14462 0 14518 800 6 la_data_in[20]
port 372 nsew signal input
rlabel metal2 s 14646 0 14702 800 6 la_data_in[21]
port 373 nsew signal input
rlabel metal2 s 14830 0 14886 800 6 la_data_in[22]
port 374 nsew signal input
rlabel metal2 s 15014 0 15070 800 6 la_data_in[23]
port 375 nsew signal input
rlabel metal2 s 15198 0 15254 800 6 la_data_in[24]
port 376 nsew signal input
rlabel metal2 s 15382 0 15438 800 6 la_data_in[25]
port 377 nsew signal input
rlabel metal2 s 15566 0 15622 800 6 la_data_in[26]
port 378 nsew signal input
rlabel metal2 s 15750 0 15806 800 6 la_data_in[27]
port 379 nsew signal input
rlabel metal2 s 15934 0 15990 800 6 la_data_in[28]
port 380 nsew signal input
rlabel metal2 s 16118 0 16174 800 6 la_data_in[29]
port 381 nsew signal input
rlabel metal2 s 11150 0 11206 800 6 la_data_in[2]
port 382 nsew signal input
rlabel metal2 s 16302 0 16358 800 6 la_data_in[30]
port 383 nsew signal input
rlabel metal2 s 16486 0 16542 800 6 la_data_in[31]
port 384 nsew signal input
rlabel metal2 s 16670 0 16726 800 6 la_data_in[32]
port 385 nsew signal input
rlabel metal2 s 16854 0 16910 800 6 la_data_in[33]
port 386 nsew signal input
rlabel metal2 s 17038 0 17094 800 6 la_data_in[34]
port 387 nsew signal input
rlabel metal2 s 17222 0 17278 800 6 la_data_in[35]
port 388 nsew signal input
rlabel metal2 s 17406 0 17462 800 6 la_data_in[36]
port 389 nsew signal input
rlabel metal2 s 17590 0 17646 800 6 la_data_in[37]
port 390 nsew signal input
rlabel metal2 s 17774 0 17830 800 6 la_data_in[38]
port 391 nsew signal input
rlabel metal2 s 17958 0 18014 800 6 la_data_in[39]
port 392 nsew signal input
rlabel metal2 s 11334 0 11390 800 6 la_data_in[3]
port 393 nsew signal input
rlabel metal2 s 18142 0 18198 800 6 la_data_in[40]
port 394 nsew signal input
rlabel metal2 s 18326 0 18382 800 6 la_data_in[41]
port 395 nsew signal input
rlabel metal2 s 18510 0 18566 800 6 la_data_in[42]
port 396 nsew signal input
rlabel metal2 s 18694 0 18750 800 6 la_data_in[43]
port 397 nsew signal input
rlabel metal2 s 18878 0 18934 800 6 la_data_in[44]
port 398 nsew signal input
rlabel metal2 s 19062 0 19118 800 6 la_data_in[45]
port 399 nsew signal input
rlabel metal2 s 19246 0 19302 800 6 la_data_in[46]
port 400 nsew signal input
rlabel metal2 s 19430 0 19486 800 6 la_data_in[47]
port 401 nsew signal input
rlabel metal2 s 19614 0 19670 800 6 la_data_in[48]
port 402 nsew signal input
rlabel metal2 s 19798 0 19854 800 6 la_data_in[49]
port 403 nsew signal input
rlabel metal2 s 11518 0 11574 800 6 la_data_in[4]
port 404 nsew signal input
rlabel metal2 s 19982 0 20038 800 6 la_data_in[50]
port 405 nsew signal input
rlabel metal2 s 20166 0 20222 800 6 la_data_in[51]
port 406 nsew signal input
rlabel metal2 s 20350 0 20406 800 6 la_data_in[52]
port 407 nsew signal input
rlabel metal2 s 20534 0 20590 800 6 la_data_in[53]
port 408 nsew signal input
rlabel metal2 s 20718 0 20774 800 6 la_data_in[54]
port 409 nsew signal input
rlabel metal2 s 20902 0 20958 800 6 la_data_in[55]
port 410 nsew signal input
rlabel metal2 s 21086 0 21142 800 6 la_data_in[56]
port 411 nsew signal input
rlabel metal2 s 21270 0 21326 800 6 la_data_in[57]
port 412 nsew signal input
rlabel metal2 s 21454 0 21510 800 6 la_data_in[58]
port 413 nsew signal input
rlabel metal2 s 21638 0 21694 800 6 la_data_in[59]
port 414 nsew signal input
rlabel metal2 s 11702 0 11758 800 6 la_data_in[5]
port 415 nsew signal input
rlabel metal2 s 21822 0 21878 800 6 la_data_in[60]
port 416 nsew signal input
rlabel metal2 s 22006 0 22062 800 6 la_data_in[61]
port 417 nsew signal input
rlabel metal2 s 22190 0 22246 800 6 la_data_in[62]
port 418 nsew signal input
rlabel metal2 s 22374 0 22430 800 6 la_data_in[63]
port 419 nsew signal input
rlabel metal2 s 22558 0 22614 800 6 la_data_in[64]
port 420 nsew signal input
rlabel metal2 s 22742 0 22798 800 6 la_data_in[65]
port 421 nsew signal input
rlabel metal2 s 22926 0 22982 800 6 la_data_in[66]
port 422 nsew signal input
rlabel metal2 s 23110 0 23166 800 6 la_data_in[67]
port 423 nsew signal input
rlabel metal2 s 23294 0 23350 800 6 la_data_in[68]
port 424 nsew signal input
rlabel metal2 s 23478 0 23534 800 6 la_data_in[69]
port 425 nsew signal input
rlabel metal2 s 11886 0 11942 800 6 la_data_in[6]
port 426 nsew signal input
rlabel metal2 s 23662 0 23718 800 6 la_data_in[70]
port 427 nsew signal input
rlabel metal2 s 23846 0 23902 800 6 la_data_in[71]
port 428 nsew signal input
rlabel metal2 s 24030 0 24086 800 6 la_data_in[72]
port 429 nsew signal input
rlabel metal2 s 24214 0 24270 800 6 la_data_in[73]
port 430 nsew signal input
rlabel metal2 s 24398 0 24454 800 6 la_data_in[74]
port 431 nsew signal input
rlabel metal2 s 24582 0 24638 800 6 la_data_in[75]
port 432 nsew signal input
rlabel metal2 s 24766 0 24822 800 6 la_data_in[76]
port 433 nsew signal input
rlabel metal2 s 24950 0 25006 800 6 la_data_in[77]
port 434 nsew signal input
rlabel metal2 s 25134 0 25190 800 6 la_data_in[78]
port 435 nsew signal input
rlabel metal2 s 25318 0 25374 800 6 la_data_in[79]
port 436 nsew signal input
rlabel metal2 s 12070 0 12126 800 6 la_data_in[7]
port 437 nsew signal input
rlabel metal2 s 25502 0 25558 800 6 la_data_in[80]
port 438 nsew signal input
rlabel metal2 s 25686 0 25742 800 6 la_data_in[81]
port 439 nsew signal input
rlabel metal2 s 25870 0 25926 800 6 la_data_in[82]
port 440 nsew signal input
rlabel metal2 s 26054 0 26110 800 6 la_data_in[83]
port 441 nsew signal input
rlabel metal2 s 26238 0 26294 800 6 la_data_in[84]
port 442 nsew signal input
rlabel metal2 s 26422 0 26478 800 6 la_data_in[85]
port 443 nsew signal input
rlabel metal2 s 26606 0 26662 800 6 la_data_in[86]
port 444 nsew signal input
rlabel metal2 s 26790 0 26846 800 6 la_data_in[87]
port 445 nsew signal input
rlabel metal2 s 26974 0 27030 800 6 la_data_in[88]
port 446 nsew signal input
rlabel metal2 s 27158 0 27214 800 6 la_data_in[89]
port 447 nsew signal input
rlabel metal2 s 12254 0 12310 800 6 la_data_in[8]
port 448 nsew signal input
rlabel metal2 s 27342 0 27398 800 6 la_data_in[90]
port 449 nsew signal input
rlabel metal2 s 27526 0 27582 800 6 la_data_in[91]
port 450 nsew signal input
rlabel metal2 s 27710 0 27766 800 6 la_data_in[92]
port 451 nsew signal input
rlabel metal2 s 27894 0 27950 800 6 la_data_in[93]
port 452 nsew signal input
rlabel metal2 s 28078 0 28134 800 6 la_data_in[94]
port 453 nsew signal input
rlabel metal2 s 28262 0 28318 800 6 la_data_in[95]
port 454 nsew signal input
rlabel metal2 s 28446 0 28502 800 6 la_data_in[96]
port 455 nsew signal input
rlabel metal2 s 28630 0 28686 800 6 la_data_in[97]
port 456 nsew signal input
rlabel metal2 s 28814 0 28870 800 6 la_data_in[98]
port 457 nsew signal input
rlabel metal2 s 28998 0 29054 800 6 la_data_in[99]
port 458 nsew signal input
rlabel metal2 s 12438 0 12494 800 6 la_data_in[9]
port 459 nsew signal input
rlabel metal2 s 34334 0 34390 800 6 la_data_out[0]
port 460 nsew signal output
rlabel metal2 s 52734 0 52790 800 6 la_data_out[100]
port 461 nsew signal output
rlabel metal2 s 52918 0 52974 800 6 la_data_out[101]
port 462 nsew signal output
rlabel metal2 s 53102 0 53158 800 6 la_data_out[102]
port 463 nsew signal output
rlabel metal2 s 53286 0 53342 800 6 la_data_out[103]
port 464 nsew signal output
rlabel metal2 s 53470 0 53526 800 6 la_data_out[104]
port 465 nsew signal output
rlabel metal2 s 53654 0 53710 800 6 la_data_out[105]
port 466 nsew signal output
rlabel metal2 s 53838 0 53894 800 6 la_data_out[106]
port 467 nsew signal output
rlabel metal2 s 54022 0 54078 800 6 la_data_out[107]
port 468 nsew signal output
rlabel metal2 s 54206 0 54262 800 6 la_data_out[108]
port 469 nsew signal output
rlabel metal2 s 54390 0 54446 800 6 la_data_out[109]
port 470 nsew signal output
rlabel metal2 s 36174 0 36230 800 6 la_data_out[10]
port 471 nsew signal output
rlabel metal2 s 54574 0 54630 800 6 la_data_out[110]
port 472 nsew signal output
rlabel metal2 s 54758 0 54814 800 6 la_data_out[111]
port 473 nsew signal output
rlabel metal2 s 54942 0 54998 800 6 la_data_out[112]
port 474 nsew signal output
rlabel metal2 s 55126 0 55182 800 6 la_data_out[113]
port 475 nsew signal output
rlabel metal2 s 55310 0 55366 800 6 la_data_out[114]
port 476 nsew signal output
rlabel metal2 s 55494 0 55550 800 6 la_data_out[115]
port 477 nsew signal output
rlabel metal2 s 55678 0 55734 800 6 la_data_out[116]
port 478 nsew signal output
rlabel metal2 s 55862 0 55918 800 6 la_data_out[117]
port 479 nsew signal output
rlabel metal2 s 56046 0 56102 800 6 la_data_out[118]
port 480 nsew signal output
rlabel metal2 s 56230 0 56286 800 6 la_data_out[119]
port 481 nsew signal output
rlabel metal2 s 36358 0 36414 800 6 la_data_out[11]
port 482 nsew signal output
rlabel metal2 s 56414 0 56470 800 6 la_data_out[120]
port 483 nsew signal output
rlabel metal2 s 56598 0 56654 800 6 la_data_out[121]
port 484 nsew signal output
rlabel metal2 s 56782 0 56838 800 6 la_data_out[122]
port 485 nsew signal output
rlabel metal2 s 56966 0 57022 800 6 la_data_out[123]
port 486 nsew signal output
rlabel metal2 s 57150 0 57206 800 6 la_data_out[124]
port 487 nsew signal output
rlabel metal2 s 57334 0 57390 800 6 la_data_out[125]
port 488 nsew signal output
rlabel metal2 s 57518 0 57574 800 6 la_data_out[126]
port 489 nsew signal output
rlabel metal2 s 57702 0 57758 800 6 la_data_out[127]
port 490 nsew signal output
rlabel metal2 s 36542 0 36598 800 6 la_data_out[12]
port 491 nsew signal output
rlabel metal2 s 36726 0 36782 800 6 la_data_out[13]
port 492 nsew signal output
rlabel metal2 s 36910 0 36966 800 6 la_data_out[14]
port 493 nsew signal output
rlabel metal2 s 37094 0 37150 800 6 la_data_out[15]
port 494 nsew signal output
rlabel metal2 s 37278 0 37334 800 6 la_data_out[16]
port 495 nsew signal output
rlabel metal2 s 37462 0 37518 800 6 la_data_out[17]
port 496 nsew signal output
rlabel metal2 s 37646 0 37702 800 6 la_data_out[18]
port 497 nsew signal output
rlabel metal2 s 37830 0 37886 800 6 la_data_out[19]
port 498 nsew signal output
rlabel metal2 s 34518 0 34574 800 6 la_data_out[1]
port 499 nsew signal output
rlabel metal2 s 38014 0 38070 800 6 la_data_out[20]
port 500 nsew signal output
rlabel metal2 s 38198 0 38254 800 6 la_data_out[21]
port 501 nsew signal output
rlabel metal2 s 38382 0 38438 800 6 la_data_out[22]
port 502 nsew signal output
rlabel metal2 s 38566 0 38622 800 6 la_data_out[23]
port 503 nsew signal output
rlabel metal2 s 38750 0 38806 800 6 la_data_out[24]
port 504 nsew signal output
rlabel metal2 s 38934 0 38990 800 6 la_data_out[25]
port 505 nsew signal output
rlabel metal2 s 39118 0 39174 800 6 la_data_out[26]
port 506 nsew signal output
rlabel metal2 s 39302 0 39358 800 6 la_data_out[27]
port 507 nsew signal output
rlabel metal2 s 39486 0 39542 800 6 la_data_out[28]
port 508 nsew signal output
rlabel metal2 s 39670 0 39726 800 6 la_data_out[29]
port 509 nsew signal output
rlabel metal2 s 34702 0 34758 800 6 la_data_out[2]
port 510 nsew signal output
rlabel metal2 s 39854 0 39910 800 6 la_data_out[30]
port 511 nsew signal output
rlabel metal2 s 40038 0 40094 800 6 la_data_out[31]
port 512 nsew signal output
rlabel metal2 s 40222 0 40278 800 6 la_data_out[32]
port 513 nsew signal output
rlabel metal2 s 40406 0 40462 800 6 la_data_out[33]
port 514 nsew signal output
rlabel metal2 s 40590 0 40646 800 6 la_data_out[34]
port 515 nsew signal output
rlabel metal2 s 40774 0 40830 800 6 la_data_out[35]
port 516 nsew signal output
rlabel metal2 s 40958 0 41014 800 6 la_data_out[36]
port 517 nsew signal output
rlabel metal2 s 41142 0 41198 800 6 la_data_out[37]
port 518 nsew signal output
rlabel metal2 s 41326 0 41382 800 6 la_data_out[38]
port 519 nsew signal output
rlabel metal2 s 41510 0 41566 800 6 la_data_out[39]
port 520 nsew signal output
rlabel metal2 s 34886 0 34942 800 6 la_data_out[3]
port 521 nsew signal output
rlabel metal2 s 41694 0 41750 800 6 la_data_out[40]
port 522 nsew signal output
rlabel metal2 s 41878 0 41934 800 6 la_data_out[41]
port 523 nsew signal output
rlabel metal2 s 42062 0 42118 800 6 la_data_out[42]
port 524 nsew signal output
rlabel metal2 s 42246 0 42302 800 6 la_data_out[43]
port 525 nsew signal output
rlabel metal2 s 42430 0 42486 800 6 la_data_out[44]
port 526 nsew signal output
rlabel metal2 s 42614 0 42670 800 6 la_data_out[45]
port 527 nsew signal output
rlabel metal2 s 42798 0 42854 800 6 la_data_out[46]
port 528 nsew signal output
rlabel metal2 s 42982 0 43038 800 6 la_data_out[47]
port 529 nsew signal output
rlabel metal2 s 43166 0 43222 800 6 la_data_out[48]
port 530 nsew signal output
rlabel metal2 s 43350 0 43406 800 6 la_data_out[49]
port 531 nsew signal output
rlabel metal2 s 35070 0 35126 800 6 la_data_out[4]
port 532 nsew signal output
rlabel metal2 s 43534 0 43590 800 6 la_data_out[50]
port 533 nsew signal output
rlabel metal2 s 43718 0 43774 800 6 la_data_out[51]
port 534 nsew signal output
rlabel metal2 s 43902 0 43958 800 6 la_data_out[52]
port 535 nsew signal output
rlabel metal2 s 44086 0 44142 800 6 la_data_out[53]
port 536 nsew signal output
rlabel metal2 s 44270 0 44326 800 6 la_data_out[54]
port 537 nsew signal output
rlabel metal2 s 44454 0 44510 800 6 la_data_out[55]
port 538 nsew signal output
rlabel metal2 s 44638 0 44694 800 6 la_data_out[56]
port 539 nsew signal output
rlabel metal2 s 44822 0 44878 800 6 la_data_out[57]
port 540 nsew signal output
rlabel metal2 s 45006 0 45062 800 6 la_data_out[58]
port 541 nsew signal output
rlabel metal2 s 45190 0 45246 800 6 la_data_out[59]
port 542 nsew signal output
rlabel metal2 s 35254 0 35310 800 6 la_data_out[5]
port 543 nsew signal output
rlabel metal2 s 45374 0 45430 800 6 la_data_out[60]
port 544 nsew signal output
rlabel metal2 s 45558 0 45614 800 6 la_data_out[61]
port 545 nsew signal output
rlabel metal2 s 45742 0 45798 800 6 la_data_out[62]
port 546 nsew signal output
rlabel metal2 s 45926 0 45982 800 6 la_data_out[63]
port 547 nsew signal output
rlabel metal2 s 46110 0 46166 800 6 la_data_out[64]
port 548 nsew signal output
rlabel metal2 s 46294 0 46350 800 6 la_data_out[65]
port 549 nsew signal output
rlabel metal2 s 46478 0 46534 800 6 la_data_out[66]
port 550 nsew signal output
rlabel metal2 s 46662 0 46718 800 6 la_data_out[67]
port 551 nsew signal output
rlabel metal2 s 46846 0 46902 800 6 la_data_out[68]
port 552 nsew signal output
rlabel metal2 s 47030 0 47086 800 6 la_data_out[69]
port 553 nsew signal output
rlabel metal2 s 35438 0 35494 800 6 la_data_out[6]
port 554 nsew signal output
rlabel metal2 s 47214 0 47270 800 6 la_data_out[70]
port 555 nsew signal output
rlabel metal2 s 47398 0 47454 800 6 la_data_out[71]
port 556 nsew signal output
rlabel metal2 s 47582 0 47638 800 6 la_data_out[72]
port 557 nsew signal output
rlabel metal2 s 47766 0 47822 800 6 la_data_out[73]
port 558 nsew signal output
rlabel metal2 s 47950 0 48006 800 6 la_data_out[74]
port 559 nsew signal output
rlabel metal2 s 48134 0 48190 800 6 la_data_out[75]
port 560 nsew signal output
rlabel metal2 s 48318 0 48374 800 6 la_data_out[76]
port 561 nsew signal output
rlabel metal2 s 48502 0 48558 800 6 la_data_out[77]
port 562 nsew signal output
rlabel metal2 s 48686 0 48742 800 6 la_data_out[78]
port 563 nsew signal output
rlabel metal2 s 48870 0 48926 800 6 la_data_out[79]
port 564 nsew signal output
rlabel metal2 s 35622 0 35678 800 6 la_data_out[7]
port 565 nsew signal output
rlabel metal2 s 49054 0 49110 800 6 la_data_out[80]
port 566 nsew signal output
rlabel metal2 s 49238 0 49294 800 6 la_data_out[81]
port 567 nsew signal output
rlabel metal2 s 49422 0 49478 800 6 la_data_out[82]
port 568 nsew signal output
rlabel metal2 s 49606 0 49662 800 6 la_data_out[83]
port 569 nsew signal output
rlabel metal2 s 49790 0 49846 800 6 la_data_out[84]
port 570 nsew signal output
rlabel metal2 s 49974 0 50030 800 6 la_data_out[85]
port 571 nsew signal output
rlabel metal2 s 50158 0 50214 800 6 la_data_out[86]
port 572 nsew signal output
rlabel metal2 s 50342 0 50398 800 6 la_data_out[87]
port 573 nsew signal output
rlabel metal2 s 50526 0 50582 800 6 la_data_out[88]
port 574 nsew signal output
rlabel metal2 s 50710 0 50766 800 6 la_data_out[89]
port 575 nsew signal output
rlabel metal2 s 35806 0 35862 800 6 la_data_out[8]
port 576 nsew signal output
rlabel metal2 s 50894 0 50950 800 6 la_data_out[90]
port 577 nsew signal output
rlabel metal2 s 51078 0 51134 800 6 la_data_out[91]
port 578 nsew signal output
rlabel metal2 s 51262 0 51318 800 6 la_data_out[92]
port 579 nsew signal output
rlabel metal2 s 51446 0 51502 800 6 la_data_out[93]
port 580 nsew signal output
rlabel metal2 s 51630 0 51686 800 6 la_data_out[94]
port 581 nsew signal output
rlabel metal2 s 51814 0 51870 800 6 la_data_out[95]
port 582 nsew signal output
rlabel metal2 s 51998 0 52054 800 6 la_data_out[96]
port 583 nsew signal output
rlabel metal2 s 52182 0 52238 800 6 la_data_out[97]
port 584 nsew signal output
rlabel metal2 s 52366 0 52422 800 6 la_data_out[98]
port 585 nsew signal output
rlabel metal2 s 52550 0 52606 800 6 la_data_out[99]
port 586 nsew signal output
rlabel metal2 s 35990 0 36046 800 6 la_data_out[9]
port 587 nsew signal output
rlabel metal3 s 67407 10072 68207 10192 6 la_oenb[0]
port 588 nsew signal input
rlabel metal3 s 0 21496 800 21616 6 la_oenb[100]
port 589 nsew signal input
rlabel metal3 s 0 22040 800 22160 6 la_oenb[101]
port 590 nsew signal input
rlabel metal3 s 0 22584 800 22704 6 la_oenb[102]
port 591 nsew signal input
rlabel metal3 s 0 23128 800 23248 6 la_oenb[103]
port 592 nsew signal input
rlabel metal3 s 0 23672 800 23792 6 la_oenb[104]
port 593 nsew signal input
rlabel metal3 s 0 24216 800 24336 6 la_oenb[105]
port 594 nsew signal input
rlabel metal3 s 0 24760 800 24880 6 la_oenb[106]
port 595 nsew signal input
rlabel metal3 s 0 25304 800 25424 6 la_oenb[107]
port 596 nsew signal input
rlabel metal3 s 0 25848 800 25968 6 la_oenb[108]
port 597 nsew signal input
rlabel metal3 s 0 26392 800 26512 6 la_oenb[109]
port 598 nsew signal input
rlabel metal3 s 67407 12792 68207 12912 6 la_oenb[10]
port 599 nsew signal input
rlabel metal3 s 0 26936 800 27056 6 la_oenb[110]
port 600 nsew signal input
rlabel metal3 s 0 27480 800 27600 6 la_oenb[111]
port 601 nsew signal input
rlabel metal3 s 0 28024 800 28144 6 la_oenb[112]
port 602 nsew signal input
rlabel metal3 s 0 28568 800 28688 6 la_oenb[113]
port 603 nsew signal input
rlabel metal3 s 0 29112 800 29232 6 la_oenb[114]
port 604 nsew signal input
rlabel metal3 s 0 29656 800 29776 6 la_oenb[115]
port 605 nsew signal input
rlabel metal3 s 0 30200 800 30320 6 la_oenb[116]
port 606 nsew signal input
rlabel metal3 s 0 30744 800 30864 6 la_oenb[117]
port 607 nsew signal input
rlabel metal3 s 0 31288 800 31408 6 la_oenb[118]
port 608 nsew signal input
rlabel metal3 s 0 31832 800 31952 6 la_oenb[119]
port 609 nsew signal input
rlabel metal3 s 67407 13064 68207 13184 6 la_oenb[11]
port 610 nsew signal input
rlabel metal3 s 0 32376 800 32496 6 la_oenb[120]
port 611 nsew signal input
rlabel metal3 s 0 32920 800 33040 6 la_oenb[121]
port 612 nsew signal input
rlabel metal3 s 0 33464 800 33584 6 la_oenb[122]
port 613 nsew signal input
rlabel metal3 s 0 34008 800 34128 6 la_oenb[123]
port 614 nsew signal input
rlabel metal3 s 0 34552 800 34672 6 la_oenb[124]
port 615 nsew signal input
rlabel metal3 s 0 35096 800 35216 6 la_oenb[125]
port 616 nsew signal input
rlabel metal3 s 0 35640 800 35760 6 la_oenb[126]
port 617 nsew signal input
rlabel metal3 s 0 36184 800 36304 6 la_oenb[127]
port 618 nsew signal input
rlabel metal3 s 67407 13336 68207 13456 6 la_oenb[12]
port 619 nsew signal input
rlabel metal3 s 67407 13608 68207 13728 6 la_oenb[13]
port 620 nsew signal input
rlabel metal3 s 67407 13880 68207 14000 6 la_oenb[14]
port 621 nsew signal input
rlabel metal3 s 67407 14152 68207 14272 6 la_oenb[15]
port 622 nsew signal input
rlabel metal3 s 67407 14424 68207 14544 6 la_oenb[16]
port 623 nsew signal input
rlabel metal3 s 67407 14696 68207 14816 6 la_oenb[17]
port 624 nsew signal input
rlabel metal3 s 67407 14968 68207 15088 6 la_oenb[18]
port 625 nsew signal input
rlabel metal3 s 67407 15240 68207 15360 6 la_oenb[19]
port 626 nsew signal input
rlabel metal3 s 67407 10344 68207 10464 6 la_oenb[1]
port 627 nsew signal input
rlabel metal3 s 67407 15512 68207 15632 6 la_oenb[20]
port 628 nsew signal input
rlabel metal3 s 67407 15784 68207 15904 6 la_oenb[21]
port 629 nsew signal input
rlabel metal3 s 67407 16056 68207 16176 6 la_oenb[22]
port 630 nsew signal input
rlabel metal3 s 67407 16328 68207 16448 6 la_oenb[23]
port 631 nsew signal input
rlabel metal3 s 67407 16600 68207 16720 6 la_oenb[24]
port 632 nsew signal input
rlabel metal3 s 67407 16872 68207 16992 6 la_oenb[25]
port 633 nsew signal input
rlabel metal3 s 67407 17144 68207 17264 6 la_oenb[26]
port 634 nsew signal input
rlabel metal3 s 67407 17416 68207 17536 6 la_oenb[27]
port 635 nsew signal input
rlabel metal3 s 67407 17688 68207 17808 6 la_oenb[28]
port 636 nsew signal input
rlabel metal3 s 67407 17960 68207 18080 6 la_oenb[29]
port 637 nsew signal input
rlabel metal3 s 67407 10616 68207 10736 6 la_oenb[2]
port 638 nsew signal input
rlabel metal3 s 67407 18232 68207 18352 6 la_oenb[30]
port 639 nsew signal input
rlabel metal3 s 67407 18504 68207 18624 6 la_oenb[31]
port 640 nsew signal input
rlabel metal3 s 67407 18776 68207 18896 6 la_oenb[32]
port 641 nsew signal input
rlabel metal3 s 67407 19048 68207 19168 6 la_oenb[33]
port 642 nsew signal input
rlabel metal3 s 67407 19320 68207 19440 6 la_oenb[34]
port 643 nsew signal input
rlabel metal3 s 67407 19592 68207 19712 6 la_oenb[35]
port 644 nsew signal input
rlabel metal3 s 67407 19864 68207 19984 6 la_oenb[36]
port 645 nsew signal input
rlabel metal3 s 67407 20136 68207 20256 6 la_oenb[37]
port 646 nsew signal input
rlabel metal3 s 67407 20408 68207 20528 6 la_oenb[38]
port 647 nsew signal input
rlabel metal3 s 67407 20680 68207 20800 6 la_oenb[39]
port 648 nsew signal input
rlabel metal3 s 67407 10888 68207 11008 6 la_oenb[3]
port 649 nsew signal input
rlabel metal3 s 67407 20952 68207 21072 6 la_oenb[40]
port 650 nsew signal input
rlabel metal3 s 67407 21224 68207 21344 6 la_oenb[41]
port 651 nsew signal input
rlabel metal3 s 67407 21496 68207 21616 6 la_oenb[42]
port 652 nsew signal input
rlabel metal3 s 67407 21768 68207 21888 6 la_oenb[43]
port 653 nsew signal input
rlabel metal3 s 67407 22040 68207 22160 6 la_oenb[44]
port 654 nsew signal input
rlabel metal3 s 67407 22312 68207 22432 6 la_oenb[45]
port 655 nsew signal input
rlabel metal3 s 67407 22584 68207 22704 6 la_oenb[46]
port 656 nsew signal input
rlabel metal3 s 67407 22856 68207 22976 6 la_oenb[47]
port 657 nsew signal input
rlabel metal3 s 67407 23128 68207 23248 6 la_oenb[48]
port 658 nsew signal input
rlabel metal3 s 67407 23400 68207 23520 6 la_oenb[49]
port 659 nsew signal input
rlabel metal3 s 67407 11160 68207 11280 6 la_oenb[4]
port 660 nsew signal input
rlabel metal3 s 67407 23672 68207 23792 6 la_oenb[50]
port 661 nsew signal input
rlabel metal3 s 67407 23944 68207 24064 6 la_oenb[51]
port 662 nsew signal input
rlabel metal3 s 67407 24216 68207 24336 6 la_oenb[52]
port 663 nsew signal input
rlabel metal3 s 67407 24488 68207 24608 6 la_oenb[53]
port 664 nsew signal input
rlabel metal3 s 67407 24760 68207 24880 6 la_oenb[54]
port 665 nsew signal input
rlabel metal3 s 67407 25032 68207 25152 6 la_oenb[55]
port 666 nsew signal input
rlabel metal3 s 67407 25304 68207 25424 6 la_oenb[56]
port 667 nsew signal input
rlabel metal3 s 67407 25576 68207 25696 6 la_oenb[57]
port 668 nsew signal input
rlabel metal3 s 67407 25848 68207 25968 6 la_oenb[58]
port 669 nsew signal input
rlabel metal3 s 67407 26120 68207 26240 6 la_oenb[59]
port 670 nsew signal input
rlabel metal3 s 67407 11432 68207 11552 6 la_oenb[5]
port 671 nsew signal input
rlabel metal3 s 67407 26392 68207 26512 6 la_oenb[60]
port 672 nsew signal input
rlabel metal3 s 67407 26664 68207 26784 6 la_oenb[61]
port 673 nsew signal input
rlabel metal3 s 67407 26936 68207 27056 6 la_oenb[62]
port 674 nsew signal input
rlabel metal3 s 67407 27208 68207 27328 6 la_oenb[63]
port 675 nsew signal input
rlabel metal3 s 67407 27480 68207 27600 6 la_oenb[64]
port 676 nsew signal input
rlabel metal3 s 67407 27752 68207 27872 6 la_oenb[65]
port 677 nsew signal input
rlabel metal3 s 67407 28024 68207 28144 6 la_oenb[66]
port 678 nsew signal input
rlabel metal3 s 67407 28296 68207 28416 6 la_oenb[67]
port 679 nsew signal input
rlabel metal3 s 67407 28568 68207 28688 6 la_oenb[68]
port 680 nsew signal input
rlabel metal3 s 0 4632 800 4752 6 la_oenb[69]
port 681 nsew signal input
rlabel metal3 s 67407 11704 68207 11824 6 la_oenb[6]
port 682 nsew signal input
rlabel metal3 s 0 5176 800 5296 6 la_oenb[70]
port 683 nsew signal input
rlabel metal3 s 0 5720 800 5840 6 la_oenb[71]
port 684 nsew signal input
rlabel metal3 s 0 6264 800 6384 6 la_oenb[72]
port 685 nsew signal input
rlabel metal3 s 0 6808 800 6928 6 la_oenb[73]
port 686 nsew signal input
rlabel metal3 s 0 7352 800 7472 6 la_oenb[74]
port 687 nsew signal input
rlabel metal3 s 0 7896 800 8016 6 la_oenb[75]
port 688 nsew signal input
rlabel metal3 s 0 8440 800 8560 6 la_oenb[76]
port 689 nsew signal input
rlabel metal3 s 0 8984 800 9104 6 la_oenb[77]
port 690 nsew signal input
rlabel metal3 s 0 9528 800 9648 6 la_oenb[78]
port 691 nsew signal input
rlabel metal3 s 0 10072 800 10192 6 la_oenb[79]
port 692 nsew signal input
rlabel metal3 s 67407 11976 68207 12096 6 la_oenb[7]
port 693 nsew signal input
rlabel metal3 s 0 10616 800 10736 6 la_oenb[80]
port 694 nsew signal input
rlabel metal3 s 0 11160 800 11280 6 la_oenb[81]
port 695 nsew signal input
rlabel metal3 s 0 11704 800 11824 6 la_oenb[82]
port 696 nsew signal input
rlabel metal3 s 0 12248 800 12368 6 la_oenb[83]
port 697 nsew signal input
rlabel metal3 s 0 12792 800 12912 6 la_oenb[84]
port 698 nsew signal input
rlabel metal3 s 0 13336 800 13456 6 la_oenb[85]
port 699 nsew signal input
rlabel metal3 s 0 13880 800 14000 6 la_oenb[86]
port 700 nsew signal input
rlabel metal3 s 0 14424 800 14544 6 la_oenb[87]
port 701 nsew signal input
rlabel metal3 s 0 14968 800 15088 6 la_oenb[88]
port 702 nsew signal input
rlabel metal3 s 0 15512 800 15632 6 la_oenb[89]
port 703 nsew signal input
rlabel metal3 s 67407 12248 68207 12368 6 la_oenb[8]
port 704 nsew signal input
rlabel metal3 s 0 16056 800 16176 6 la_oenb[90]
port 705 nsew signal input
rlabel metal3 s 0 16600 800 16720 6 la_oenb[91]
port 706 nsew signal input
rlabel metal3 s 0 17144 800 17264 6 la_oenb[92]
port 707 nsew signal input
rlabel metal3 s 0 17688 800 17808 6 la_oenb[93]
port 708 nsew signal input
rlabel metal3 s 0 18232 800 18352 6 la_oenb[94]
port 709 nsew signal input
rlabel metal3 s 0 18776 800 18896 6 la_oenb[95]
port 710 nsew signal input
rlabel metal3 s 0 19320 800 19440 6 la_oenb[96]
port 711 nsew signal input
rlabel metal3 s 0 19864 800 19984 6 la_oenb[97]
port 712 nsew signal input
rlabel metal3 s 0 20408 800 20528 6 la_oenb[98]
port 713 nsew signal input
rlabel metal3 s 0 20952 800 21072 6 la_oenb[99]
port 714 nsew signal input
rlabel metal3 s 67407 12520 68207 12640 6 la_oenb[9]
port 715 nsew signal input
rlabel metal3 s 0 1368 800 1488 6 load_data
port 716 nsew signal output
rlabel metal3 s 0 3000 800 3120 6 load_status[0]
port 717 nsew signal output
rlabel metal3 s 0 3544 800 3664 6 load_status[1]
port 718 nsew signal output
rlabel metal3 s 0 4088 800 4208 6 load_status[2]
port 719 nsew signal output
rlabel metal3 s 0 824 800 944 6 master_ena_proc
port 720 nsew signal output
rlabel metal3 s 67407 8712 68207 8832 6 next_key
port 721 nsew signal input
rlabel metal3 s 67407 8440 68207 8560 6 slv_done
port 722 nsew signal input
rlabel metal3 s 0 1912 800 2032 6 trigLoad
port 723 nsew signal output
rlabel metal4 s 9189 2128 9509 34864 6 vccd1
port 724 nsew power bidirectional
rlabel metal4 s 25680 2128 26000 34864 6 vccd1
port 724 nsew power bidirectional
rlabel metal4 s 42171 2128 42491 34864 6 vccd1
port 724 nsew power bidirectional
rlabel metal4 s 58662 2128 58982 34864 6 vccd1
port 724 nsew power bidirectional
rlabel metal4 s 17434 2128 17754 34864 6 vssd1
port 725 nsew ground bidirectional
rlabel metal4 s 33925 2128 34245 34864 6 vssd1
port 725 nsew ground bidirectional
rlabel metal4 s 50416 2128 50736 34864 6 vssd1
port 725 nsew ground bidirectional
rlabel metal4 s 66907 2128 67227 34864 6 vssd1
port 725 nsew ground bidirectional
rlabel metal2 s 10414 0 10470 800 6 wb_clk_i
port 726 nsew signal input
rlabel metal2 s 10598 0 10654 800 6 wb_rst_i
port 727 nsew signal input
<< properties >>
string FIXED_BBOX 0 0 68207 37351
string LEFclass BLOCK
string LEFview TRUE
string GDS_END 9656726
string GDS_FILE /mnt/d/BEC/bec-unic/openlane/controller/runs/24_10_20_04_20/results/signoff/controller.magic.gds
string GDS_START 547748
<< end >>

