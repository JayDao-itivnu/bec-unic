// This is the unpowered netlist.
module controller (ki,
    load_data,
    master_ena_proc,
    next_key,
    slv_done,
    trigLoad,
    wb_clk_i,
    wb_rst_i,
    becStatus,
    data_in,
    data_out,
    la_data_in,
    la_data_out,
    la_oenb,
    load_status);
 output ki;
 output load_data;
 output master_ena_proc;
 input next_key;
 input slv_done;
 output trigLoad;
 input wb_clk_i;
 input wb_rst_i;
 input [3:0] becStatus;
 input [162:0] data_in;
 output [162:0] data_out;
 input [127:0] la_data_in;
 output [127:0] la_data_out;
 input [127:0] la_oenb;
 output [2:0] load_status;

 wire net618;
 wire net628;
 wire net650;
 wire net651;
 wire net652;
 wire net653;
 wire net654;
 wire net655;
 wire net629;
 wire net656;
 wire net657;
 wire net630;
 wire net631;
 wire net632;
 wire net633;
 wire net634;
 wire net635;
 wire net636;
 wire net637;
 wire net619;
 wire net638;
 wire net639;
 wire net640;
 wire net641;
 wire net642;
 wire net643;
 wire net644;
 wire net645;
 wire net646;
 wire net647;
 wire net620;
 wire net648;
 wire net649;
 wire net621;
 wire net622;
 wire net623;
 wire net624;
 wire net625;
 wire net626;
 wire net627;
 wire _0000_;
 wire _0001_;
 wire _0002_;
 wire _0003_;
 wire _0004_;
 wire _0005_;
 wire _0006_;
 wire _0007_;
 wire _0008_;
 wire _0009_;
 wire _0010_;
 wire _0011_;
 wire _0012_;
 wire _0013_;
 wire _0014_;
 wire _0015_;
 wire _0016_;
 wire _0017_;
 wire _0018_;
 wire _0019_;
 wire _0020_;
 wire _0021_;
 wire _0022_;
 wire _0023_;
 wire _0024_;
 wire _0025_;
 wire _0026_;
 wire _0027_;
 wire _0028_;
 wire _0029_;
 wire _0030_;
 wire _0031_;
 wire _0032_;
 wire _0033_;
 wire _0034_;
 wire _0035_;
 wire _0036_;
 wire _0037_;
 wire _0038_;
 wire _0039_;
 wire _0040_;
 wire _0041_;
 wire _0042_;
 wire _0043_;
 wire _0044_;
 wire _0045_;
 wire _0046_;
 wire _0047_;
 wire _0048_;
 wire _0049_;
 wire _0050_;
 wire _0051_;
 wire _0052_;
 wire _0053_;
 wire _0054_;
 wire _0055_;
 wire _0056_;
 wire _0057_;
 wire _0058_;
 wire _0059_;
 wire _0060_;
 wire _0061_;
 wire _0062_;
 wire _0063_;
 wire _0064_;
 wire _0065_;
 wire _0066_;
 wire _0067_;
 wire _0068_;
 wire _0069_;
 wire _0070_;
 wire _0071_;
 wire _0072_;
 wire _0073_;
 wire _0074_;
 wire _0075_;
 wire _0076_;
 wire _0077_;
 wire _0078_;
 wire _0079_;
 wire _0080_;
 wire _0081_;
 wire _0082_;
 wire _0083_;
 wire _0084_;
 wire _0085_;
 wire _0086_;
 wire _0087_;
 wire _0088_;
 wire _0089_;
 wire _0090_;
 wire _0091_;
 wire _0092_;
 wire _0093_;
 wire _0094_;
 wire _0095_;
 wire _0096_;
 wire _0097_;
 wire _0098_;
 wire _0099_;
 wire _0100_;
 wire _0101_;
 wire _0102_;
 wire _0103_;
 wire _0104_;
 wire _0105_;
 wire _0106_;
 wire _0107_;
 wire _0108_;
 wire _0109_;
 wire _0110_;
 wire _0111_;
 wire _0112_;
 wire _0113_;
 wire _0114_;
 wire _0115_;
 wire _0116_;
 wire _0117_;
 wire _0118_;
 wire _0119_;
 wire _0120_;
 wire _0121_;
 wire _0122_;
 wire _0123_;
 wire _0124_;
 wire _0125_;
 wire _0126_;
 wire _0127_;
 wire _0128_;
 wire _0129_;
 wire _0130_;
 wire _0131_;
 wire _0132_;
 wire _0133_;
 wire _0134_;
 wire _0135_;
 wire _0136_;
 wire _0137_;
 wire _0138_;
 wire _0139_;
 wire _0140_;
 wire _0141_;
 wire _0142_;
 wire _0143_;
 wire _0144_;
 wire _0145_;
 wire _0146_;
 wire _0147_;
 wire _0148_;
 wire _0149_;
 wire _0150_;
 wire _0151_;
 wire _0152_;
 wire _0153_;
 wire _0154_;
 wire _0155_;
 wire _0156_;
 wire _0157_;
 wire _0158_;
 wire _0159_;
 wire _0160_;
 wire _0161_;
 wire _0162_;
 wire _0163_;
 wire _0164_;
 wire _0165_;
 wire _0166_;
 wire _0167_;
 wire _0168_;
 wire _0169_;
 wire _0170_;
 wire _0171_;
 wire _0172_;
 wire _0173_;
 wire _0174_;
 wire _0175_;
 wire _0176_;
 wire _0177_;
 wire _0178_;
 wire _0179_;
 wire _0180_;
 wire _0181_;
 wire _0182_;
 wire _0183_;
 wire _0184_;
 wire _0185_;
 wire _0186_;
 wire _0187_;
 wire _0188_;
 wire _0189_;
 wire _0190_;
 wire _0191_;
 wire _0192_;
 wire _0193_;
 wire _0194_;
 wire _0195_;
 wire _0196_;
 wire _0197_;
 wire _0198_;
 wire _0199_;
 wire _0200_;
 wire _0201_;
 wire _0202_;
 wire _0203_;
 wire _0204_;
 wire _0205_;
 wire _0206_;
 wire _0207_;
 wire _0208_;
 wire _0209_;
 wire _0210_;
 wire _0211_;
 wire _0212_;
 wire _0213_;
 wire _0214_;
 wire _0215_;
 wire _0216_;
 wire _0217_;
 wire _0218_;
 wire _0219_;
 wire _0220_;
 wire _0221_;
 wire _0222_;
 wire _0223_;
 wire _0224_;
 wire _0225_;
 wire _0226_;
 wire _0227_;
 wire _0228_;
 wire _0229_;
 wire _0230_;
 wire _0231_;
 wire _0232_;
 wire _0233_;
 wire _0234_;
 wire _0235_;
 wire _0236_;
 wire _0237_;
 wire _0238_;
 wire _0239_;
 wire _0240_;
 wire _0241_;
 wire _0242_;
 wire _0243_;
 wire _0244_;
 wire _0245_;
 wire _0246_;
 wire _0247_;
 wire _0248_;
 wire _0249_;
 wire _0250_;
 wire _0251_;
 wire _0252_;
 wire _0253_;
 wire _0254_;
 wire _0255_;
 wire _0256_;
 wire _0257_;
 wire _0258_;
 wire _0259_;
 wire _0260_;
 wire _0261_;
 wire _0262_;
 wire _0263_;
 wire _0264_;
 wire _0265_;
 wire _0266_;
 wire _0267_;
 wire _0268_;
 wire _0269_;
 wire _0270_;
 wire _0271_;
 wire _0272_;
 wire _0273_;
 wire _0274_;
 wire _0275_;
 wire _0276_;
 wire _0277_;
 wire _0278_;
 wire _0279_;
 wire _0280_;
 wire _0281_;
 wire _0282_;
 wire _0283_;
 wire _0284_;
 wire _0285_;
 wire _0286_;
 wire _0287_;
 wire _0288_;
 wire _0289_;
 wire _0290_;
 wire _0291_;
 wire _0292_;
 wire _0293_;
 wire _0294_;
 wire _0295_;
 wire _0296_;
 wire _0297_;
 wire _0298_;
 wire _0299_;
 wire _0300_;
 wire _0301_;
 wire _0302_;
 wire _0303_;
 wire _0304_;
 wire _0305_;
 wire _0306_;
 wire _0307_;
 wire _0308_;
 wire _0309_;
 wire _0310_;
 wire _0311_;
 wire _0312_;
 wire _0313_;
 wire _0314_;
 wire _0315_;
 wire _0316_;
 wire _0317_;
 wire _0318_;
 wire _0319_;
 wire _0320_;
 wire _0321_;
 wire _0322_;
 wire _0323_;
 wire _0324_;
 wire _0325_;
 wire _0326_;
 wire _0327_;
 wire _0328_;
 wire _0329_;
 wire _0330_;
 wire _0331_;
 wire _0332_;
 wire _0333_;
 wire _0334_;
 wire _0335_;
 wire _0336_;
 wire _0337_;
 wire _0338_;
 wire _0339_;
 wire _0340_;
 wire _0341_;
 wire _0342_;
 wire _0343_;
 wire _0344_;
 wire _0345_;
 wire _0346_;
 wire _0347_;
 wire _0348_;
 wire _0349_;
 wire _0350_;
 wire _0351_;
 wire _0352_;
 wire _0353_;
 wire _0354_;
 wire _0355_;
 wire _0356_;
 wire _0357_;
 wire _0358_;
 wire _0359_;
 wire _0360_;
 wire _0361_;
 wire _0362_;
 wire _0363_;
 wire _0364_;
 wire _0365_;
 wire _0366_;
 wire _0367_;
 wire _0368_;
 wire _0369_;
 wire _0370_;
 wire _0371_;
 wire _0372_;
 wire _0373_;
 wire _0374_;
 wire _0375_;
 wire _0376_;
 wire _0377_;
 wire _0378_;
 wire _0379_;
 wire _0380_;
 wire _0381_;
 wire _0382_;
 wire _0383_;
 wire _0384_;
 wire _0385_;
 wire _0386_;
 wire _0387_;
 wire _0388_;
 wire _0389_;
 wire _0390_;
 wire _0391_;
 wire _0392_;
 wire _0393_;
 wire _0394_;
 wire _0395_;
 wire _0396_;
 wire _0397_;
 wire _0398_;
 wire _0399_;
 wire _0400_;
 wire _0401_;
 wire _0402_;
 wire _0403_;
 wire _0404_;
 wire _0405_;
 wire _0406_;
 wire _0407_;
 wire _0408_;
 wire _0409_;
 wire _0410_;
 wire _0411_;
 wire _0412_;
 wire _0413_;
 wire _0414_;
 wire _0415_;
 wire _0416_;
 wire _0417_;
 wire _0418_;
 wire _0419_;
 wire _0420_;
 wire _0421_;
 wire _0422_;
 wire _0423_;
 wire _0424_;
 wire _0425_;
 wire _0426_;
 wire _0427_;
 wire _0428_;
 wire _0429_;
 wire _0430_;
 wire _0431_;
 wire _0432_;
 wire _0433_;
 wire _0434_;
 wire _0435_;
 wire _0436_;
 wire _0437_;
 wire _0438_;
 wire _0439_;
 wire _0440_;
 wire _0441_;
 wire _0442_;
 wire _0443_;
 wire _0444_;
 wire _0445_;
 wire _0446_;
 wire _0447_;
 wire _0448_;
 wire _0449_;
 wire _0450_;
 wire _0451_;
 wire _0452_;
 wire _0453_;
 wire _0454_;
 wire _0455_;
 wire _0456_;
 wire _0457_;
 wire _0458_;
 wire _0459_;
 wire _0460_;
 wire _0461_;
 wire _0462_;
 wire _0463_;
 wire _0464_;
 wire _0465_;
 wire _0466_;
 wire _0467_;
 wire _0468_;
 wire _0469_;
 wire _0470_;
 wire _0471_;
 wire _0472_;
 wire _0473_;
 wire _0474_;
 wire _0475_;
 wire _0476_;
 wire _0477_;
 wire _0478_;
 wire _0479_;
 wire _0480_;
 wire _0481_;
 wire _0482_;
 wire _0483_;
 wire _0484_;
 wire _0485_;
 wire _0486_;
 wire _0487_;
 wire _0488_;
 wire _0489_;
 wire _0490_;
 wire _0491_;
 wire _0492_;
 wire _0493_;
 wire _0494_;
 wire _0495_;
 wire _0496_;
 wire _0497_;
 wire _0498_;
 wire _0499_;
 wire _0500_;
 wire _0501_;
 wire _0502_;
 wire _0503_;
 wire _0504_;
 wire _0505_;
 wire _0506_;
 wire _0507_;
 wire _0508_;
 wire _0509_;
 wire _0510_;
 wire _0511_;
 wire _0512_;
 wire _0513_;
 wire _0514_;
 wire _0515_;
 wire _0516_;
 wire _0517_;
 wire _0518_;
 wire _0519_;
 wire _0520_;
 wire _0521_;
 wire _0522_;
 wire _0523_;
 wire _0524_;
 wire _0525_;
 wire _0526_;
 wire _0527_;
 wire _0528_;
 wire _0529_;
 wire _0530_;
 wire _0531_;
 wire _0532_;
 wire _0533_;
 wire _0534_;
 wire _0535_;
 wire _0536_;
 wire _0537_;
 wire _0538_;
 wire _0539_;
 wire _0540_;
 wire _0541_;
 wire _0542_;
 wire _0543_;
 wire _0544_;
 wire _0545_;
 wire _0546_;
 wire _0547_;
 wire _0548_;
 wire _0549_;
 wire _0550_;
 wire _0551_;
 wire _0552_;
 wire _0553_;
 wire _0554_;
 wire _0555_;
 wire _0556_;
 wire _0557_;
 wire _0558_;
 wire _0559_;
 wire _0560_;
 wire _0561_;
 wire _0562_;
 wire _0563_;
 wire _0564_;
 wire _0565_;
 wire _0566_;
 wire _0567_;
 wire _0568_;
 wire _0569_;
 wire _0570_;
 wire _0571_;
 wire _0572_;
 wire _0573_;
 wire _0574_;
 wire _0575_;
 wire _0576_;
 wire _0577_;
 wire _0578_;
 wire _0579_;
 wire _0580_;
 wire _0581_;
 wire _0582_;
 wire _0583_;
 wire _0584_;
 wire _0585_;
 wire _0586_;
 wire _0587_;
 wire _0588_;
 wire _0589_;
 wire _0590_;
 wire _0591_;
 wire _0592_;
 wire _0593_;
 wire _0594_;
 wire _0595_;
 wire _0596_;
 wire _0597_;
 wire _0598_;
 wire _0599_;
 wire _0600_;
 wire _0601_;
 wire _0602_;
 wire _0603_;
 wire _0604_;
 wire _0605_;
 wire _0606_;
 wire _0607_;
 wire _0608_;
 wire _0609_;
 wire _0610_;
 wire _0611_;
 wire _0612_;
 wire _0613_;
 wire _0614_;
 wire _0615_;
 wire _0616_;
 wire _0617_;
 wire _0618_;
 wire _0619_;
 wire _0620_;
 wire _0621_;
 wire _0622_;
 wire _0623_;
 wire _0624_;
 wire _0625_;
 wire _0626_;
 wire _0627_;
 wire _0628_;
 wire _0629_;
 wire _0630_;
 wire _0631_;
 wire _0632_;
 wire _0633_;
 wire _0634_;
 wire _0635_;
 wire _0636_;
 wire _0637_;
 wire _0638_;
 wire _0639_;
 wire _0640_;
 wire _0641_;
 wire _0642_;
 wire _0643_;
 wire _0644_;
 wire _0645_;
 wire _0646_;
 wire _0647_;
 wire _0648_;
 wire _0649_;
 wire _0650_;
 wire _0651_;
 wire _0652_;
 wire _0653_;
 wire _0654_;
 wire _0655_;
 wire _0656_;
 wire _0657_;
 wire _0658_;
 wire _0659_;
 wire _0660_;
 wire _0661_;
 wire _0662_;
 wire _0663_;
 wire _0664_;
 wire _0665_;
 wire _0666_;
 wire _0667_;
 wire _0668_;
 wire _0669_;
 wire _0670_;
 wire _0671_;
 wire _0672_;
 wire _0673_;
 wire _0674_;
 wire _0675_;
 wire _0676_;
 wire _0677_;
 wire _0678_;
 wire _0679_;
 wire _0680_;
 wire _0681_;
 wire _0682_;
 wire _0683_;
 wire _0684_;
 wire _0685_;
 wire _0686_;
 wire _0687_;
 wire _0688_;
 wire _0689_;
 wire _0690_;
 wire _0691_;
 wire _0692_;
 wire _0693_;
 wire _0694_;
 wire _0695_;
 wire _0696_;
 wire _0697_;
 wire _0698_;
 wire _0699_;
 wire _0700_;
 wire _0701_;
 wire _0702_;
 wire _0703_;
 wire _0704_;
 wire _0705_;
 wire _0706_;
 wire _0707_;
 wire _0708_;
 wire _0709_;
 wire _0710_;
 wire _0711_;
 wire _0712_;
 wire _0713_;
 wire _0714_;
 wire _0715_;
 wire _0716_;
 wire _0717_;
 wire _0718_;
 wire _0719_;
 wire _0720_;
 wire _0721_;
 wire _0722_;
 wire _0723_;
 wire _0724_;
 wire _0725_;
 wire _0726_;
 wire _0727_;
 wire _0728_;
 wire _0729_;
 wire _0730_;
 wire _0731_;
 wire _0732_;
 wire _0733_;
 wire _0734_;
 wire _0735_;
 wire _0736_;
 wire _0737_;
 wire _0738_;
 wire _0739_;
 wire _0740_;
 wire _0741_;
 wire _0742_;
 wire _0743_;
 wire _0744_;
 wire _0745_;
 wire _0746_;
 wire _0747_;
 wire _0748_;
 wire _0749_;
 wire _0750_;
 wire _0751_;
 wire _0752_;
 wire _0753_;
 wire _0754_;
 wire _0755_;
 wire _0756_;
 wire _0757_;
 wire _0758_;
 wire _0759_;
 wire _0760_;
 wire _0761_;
 wire _0762_;
 wire _0763_;
 wire _0764_;
 wire _0765_;
 wire _0766_;
 wire _0767_;
 wire _0768_;
 wire _0769_;
 wire _0770_;
 wire _0771_;
 wire _0772_;
 wire _0773_;
 wire _0774_;
 wire _0775_;
 wire _0776_;
 wire _0777_;
 wire _0778_;
 wire _0779_;
 wire _0780_;
 wire _0781_;
 wire _0782_;
 wire _0783_;
 wire _0784_;
 wire _0785_;
 wire _0786_;
 wire _0787_;
 wire _0788_;
 wire _0789_;
 wire _0790_;
 wire _0791_;
 wire _0792_;
 wire _0793_;
 wire _0794_;
 wire _0795_;
 wire _0796_;
 wire _0797_;
 wire _0798_;
 wire _0799_;
 wire _0800_;
 wire _0801_;
 wire _0802_;
 wire _0803_;
 wire _0804_;
 wire _0805_;
 wire _0806_;
 wire _0807_;
 wire _0808_;
 wire _0809_;
 wire _0810_;
 wire _0811_;
 wire _0812_;
 wire _0813_;
 wire _0814_;
 wire _0815_;
 wire _0816_;
 wire _0817_;
 wire _0818_;
 wire _0819_;
 wire _0820_;
 wire _0821_;
 wire _0822_;
 wire _0823_;
 wire _0824_;
 wire _0825_;
 wire _0826_;
 wire _0827_;
 wire _0828_;
 wire _0829_;
 wire _0830_;
 wire _0831_;
 wire _0832_;
 wire _0833_;
 wire _0834_;
 wire _0835_;
 wire _0836_;
 wire _0837_;
 wire _0838_;
 wire _0839_;
 wire _0840_;
 wire _0841_;
 wire _0842_;
 wire _0843_;
 wire _0844_;
 wire _0845_;
 wire _0846_;
 wire _0847_;
 wire _0848_;
 wire _0849_;
 wire _0850_;
 wire _0851_;
 wire _0852_;
 wire _0853_;
 wire _0854_;
 wire _0855_;
 wire _0856_;
 wire _0857_;
 wire _0858_;
 wire _0859_;
 wire _0860_;
 wire _0861_;
 wire _0862_;
 wire _0863_;
 wire _0864_;
 wire _0865_;
 wire _0866_;
 wire _0867_;
 wire _0868_;
 wire _0869_;
 wire _0870_;
 wire _0871_;
 wire _0872_;
 wire _0873_;
 wire _0874_;
 wire _0875_;
 wire _0876_;
 wire _0877_;
 wire _0878_;
 wire _0879_;
 wire _0880_;
 wire _0881_;
 wire _0882_;
 wire _0883_;
 wire _0884_;
 wire _0885_;
 wire _0886_;
 wire _0887_;
 wire _0888_;
 wire _0889_;
 wire _0890_;
 wire _0891_;
 wire _0892_;
 wire _0893_;
 wire _0894_;
 wire _0895_;
 wire _0896_;
 wire _0897_;
 wire _0898_;
 wire _0899_;
 wire _0900_;
 wire _0901_;
 wire _0902_;
 wire _0903_;
 wire _0904_;
 wire _0905_;
 wire _0906_;
 wire _0907_;
 wire _0908_;
 wire _0909_;
 wire _0910_;
 wire _0911_;
 wire _0912_;
 wire _0913_;
 wire _0914_;
 wire _0915_;
 wire _0916_;
 wire _0917_;
 wire _0918_;
 wire _0919_;
 wire _0920_;
 wire _0921_;
 wire _0922_;
 wire _0923_;
 wire _0924_;
 wire _0925_;
 wire _0926_;
 wire _0927_;
 wire _0928_;
 wire _0929_;
 wire _0930_;
 wire _0931_;
 wire _0932_;
 wire _0933_;
 wire _0934_;
 wire _0935_;
 wire _0936_;
 wire _0937_;
 wire _0938_;
 wire _0939_;
 wire _0940_;
 wire _0941_;
 wire _0942_;
 wire _0943_;
 wire _0944_;
 wire _0945_;
 wire _0946_;
 wire _0947_;
 wire _0948_;
 wire _0949_;
 wire _0950_;
 wire _0951_;
 wire clknet_0_wb_clk_i;
 wire clknet_1_0__leaf_wb_clk_i;
 wire clknet_1_1__leaf_wb_clk_i;
 wire clknet_leaf_0_wb_clk_i;
 wire clknet_leaf_10_wb_clk_i;
 wire clknet_leaf_11_wb_clk_i;
 wire clknet_leaf_12_wb_clk_i;
 wire clknet_leaf_13_wb_clk_i;
 wire clknet_leaf_14_wb_clk_i;
 wire clknet_leaf_15_wb_clk_i;
 wire clknet_leaf_16_wb_clk_i;
 wire clknet_leaf_17_wb_clk_i;
 wire clknet_leaf_18_wb_clk_i;
 wire clknet_leaf_19_wb_clk_i;
 wire clknet_leaf_1_wb_clk_i;
 wire clknet_leaf_20_wb_clk_i;
 wire clknet_leaf_21_wb_clk_i;
 wire clknet_leaf_22_wb_clk_i;
 wire clknet_leaf_23_wb_clk_i;
 wire clknet_leaf_24_wb_clk_i;
 wire clknet_leaf_25_wb_clk_i;
 wire clknet_leaf_26_wb_clk_i;
 wire clknet_leaf_2_wb_clk_i;
 wire clknet_leaf_3_wb_clk_i;
 wire clknet_leaf_4_wb_clk_i;
 wire clknet_leaf_5_wb_clk_i;
 wire clknet_leaf_6_wb_clk_i;
 wire clknet_leaf_7_wb_clk_i;
 wire clknet_leaf_8_wb_clk_i;
 wire clknet_leaf_9_wb_clk_i;
 wire \current_state[0] ;
 wire \current_state[1] ;
 wire enable_proc;
 wire net1;
 wire net10;
 wire net100;
 wire net1000;
 wire net1001;
 wire net1002;
 wire net1003;
 wire net1004;
 wire net1005;
 wire net1006;
 wire net1007;
 wire net1008;
 wire net1009;
 wire net101;
 wire net1010;
 wire net1011;
 wire net1012;
 wire net1013;
 wire net1014;
 wire net1015;
 wire net1016;
 wire net1017;
 wire net1018;
 wire net1019;
 wire net102;
 wire net1020;
 wire net1021;
 wire net1022;
 wire net1023;
 wire net1024;
 wire net1025;
 wire net1026;
 wire net1027;
 wire net1028;
 wire net1029;
 wire net103;
 wire net1030;
 wire net1031;
 wire net1032;
 wire net1033;
 wire net1034;
 wire net1035;
 wire net1036;
 wire net1037;
 wire net1038;
 wire net1039;
 wire net104;
 wire net1040;
 wire net1041;
 wire net1042;
 wire net1043;
 wire net1044;
 wire net1045;
 wire net1046;
 wire net1047;
 wire net1048;
 wire net1049;
 wire net105;
 wire net1050;
 wire net1051;
 wire net1052;
 wire net1053;
 wire net1054;
 wire net1055;
 wire net1056;
 wire net1057;
 wire net1058;
 wire net1059;
 wire net106;
 wire net1060;
 wire net1061;
 wire net1062;
 wire net1063;
 wire net1064;
 wire net1065;
 wire net1066;
 wire net1067;
 wire net1068;
 wire net1069;
 wire net107;
 wire net1070;
 wire net1071;
 wire net1072;
 wire net1073;
 wire net1074;
 wire net1075;
 wire net1076;
 wire net1077;
 wire net1078;
 wire net1079;
 wire net108;
 wire net1080;
 wire net1081;
 wire net1082;
 wire net1083;
 wire net1084;
 wire net1085;
 wire net1086;
 wire net1087;
 wire net1088;
 wire net1089;
 wire net109;
 wire net1090;
 wire net1091;
 wire net1092;
 wire net1093;
 wire net1094;
 wire net1095;
 wire net1096;
 wire net1097;
 wire net1098;
 wire net1099;
 wire net11;
 wire net110;
 wire net1100;
 wire net1101;
 wire net1102;
 wire net1103;
 wire net1104;
 wire net1105;
 wire net1106;
 wire net1107;
 wire net1108;
 wire net1109;
 wire net111;
 wire net1110;
 wire net1111;
 wire net1112;
 wire net1113;
 wire net1114;
 wire net1115;
 wire net1116;
 wire net1117;
 wire net1118;
 wire net1119;
 wire net112;
 wire net1120;
 wire net1121;
 wire net1122;
 wire net1123;
 wire net1124;
 wire net1125;
 wire net1126;
 wire net1127;
 wire net1128;
 wire net1129;
 wire net113;
 wire net1130;
 wire net1131;
 wire net1132;
 wire net1133;
 wire net1134;
 wire net1135;
 wire net1136;
 wire net1137;
 wire net1138;
 wire net1139;
 wire net114;
 wire net1140;
 wire net1141;
 wire net1142;
 wire net1143;
 wire net1144;
 wire net1145;
 wire net1146;
 wire net1147;
 wire net1148;
 wire net1149;
 wire net115;
 wire net1150;
 wire net1151;
 wire net1152;
 wire net1153;
 wire net1154;
 wire net1155;
 wire net1156;
 wire net1157;
 wire net1158;
 wire net1159;
 wire net116;
 wire net1160;
 wire net1161;
 wire net1162;
 wire net1163;
 wire net1164;
 wire net1165;
 wire net1166;
 wire net1167;
 wire net1168;
 wire net1169;
 wire net117;
 wire net1170;
 wire net1171;
 wire net1172;
 wire net1173;
 wire net1174;
 wire net1175;
 wire net1176;
 wire net1177;
 wire net1178;
 wire net1179;
 wire net118;
 wire net1180;
 wire net1181;
 wire net1182;
 wire net1183;
 wire net1184;
 wire net1185;
 wire net1186;
 wire net1187;
 wire net1188;
 wire net1189;
 wire net119;
 wire net1190;
 wire net1191;
 wire net1192;
 wire net1193;
 wire net1194;
 wire net1195;
 wire net1196;
 wire net1197;
 wire net1198;
 wire net1199;
 wire net12;
 wire net120;
 wire net1200;
 wire net1201;
 wire net1202;
 wire net1203;
 wire net1204;
 wire net1205;
 wire net1206;
 wire net1207;
 wire net1208;
 wire net1209;
 wire net121;
 wire net1210;
 wire net1211;
 wire net1212;
 wire net1213;
 wire net1214;
 wire net1215;
 wire net1216;
 wire net1217;
 wire net1218;
 wire net1219;
 wire net122;
 wire net1220;
 wire net1221;
 wire net1222;
 wire net1223;
 wire net1224;
 wire net1225;
 wire net1226;
 wire net1227;
 wire net1228;
 wire net1229;
 wire net123;
 wire net1230;
 wire net1231;
 wire net1232;
 wire net1233;
 wire net1234;
 wire net1235;
 wire net1236;
 wire net1237;
 wire net1238;
 wire net1239;
 wire net124;
 wire net1240;
 wire net1241;
 wire net1242;
 wire net1243;
 wire net1244;
 wire net1245;
 wire net1246;
 wire net1247;
 wire net1248;
 wire net1249;
 wire net125;
 wire net1250;
 wire net1251;
 wire net1252;
 wire net1253;
 wire net1254;
 wire net1255;
 wire net1256;
 wire net1257;
 wire net1258;
 wire net1259;
 wire net126;
 wire net1260;
 wire net1261;
 wire net1262;
 wire net1263;
 wire net1264;
 wire net1265;
 wire net1266;
 wire net1267;
 wire net1268;
 wire net1269;
 wire net127;
 wire net1270;
 wire net1271;
 wire net1272;
 wire net1273;
 wire net1274;
 wire net1275;
 wire net1276;
 wire net1277;
 wire net1278;
 wire net1279;
 wire net128;
 wire net1280;
 wire net1281;
 wire net1282;
 wire net1283;
 wire net1284;
 wire net1285;
 wire net1286;
 wire net1287;
 wire net1288;
 wire net1289;
 wire net129;
 wire net1290;
 wire net1291;
 wire net1292;
 wire net1293;
 wire net1294;
 wire net1295;
 wire net1296;
 wire net1297;
 wire net1298;
 wire net1299;
 wire net13;
 wire net130;
 wire net1300;
 wire net1301;
 wire net1302;
 wire net1303;
 wire net1304;
 wire net1305;
 wire net1306;
 wire net1307;
 wire net1308;
 wire net1309;
 wire net131;
 wire net1310;
 wire net1311;
 wire net1312;
 wire net1313;
 wire net1314;
 wire net1315;
 wire net1316;
 wire net1317;
 wire net1318;
 wire net1319;
 wire net132;
 wire net1320;
 wire net1321;
 wire net1322;
 wire net1323;
 wire net1324;
 wire net1325;
 wire net1326;
 wire net1327;
 wire net1328;
 wire net1329;
 wire net133;
 wire net1330;
 wire net1331;
 wire net1332;
 wire net1333;
 wire net1334;
 wire net1335;
 wire net1336;
 wire net1337;
 wire net1338;
 wire net1339;
 wire net134;
 wire net1340;
 wire net1341;
 wire net1342;
 wire net1343;
 wire net1344;
 wire net1345;
 wire net1346;
 wire net1347;
 wire net1348;
 wire net1349;
 wire net135;
 wire net1350;
 wire net1351;
 wire net1352;
 wire net1353;
 wire net1354;
 wire net1355;
 wire net1356;
 wire net1357;
 wire net1358;
 wire net1359;
 wire net136;
 wire net1360;
 wire net1361;
 wire net1362;
 wire net1363;
 wire net1364;
 wire net1365;
 wire net1366;
 wire net1367;
 wire net1368;
 wire net1369;
 wire net137;
 wire net1370;
 wire net1371;
 wire net1372;
 wire net1373;
 wire net1374;
 wire net1375;
 wire net1376;
 wire net1377;
 wire net1378;
 wire net1379;
 wire net138;
 wire net1380;
 wire net1381;
 wire net1382;
 wire net1383;
 wire net1384;
 wire net1385;
 wire net1386;
 wire net1387;
 wire net1388;
 wire net1389;
 wire net139;
 wire net1390;
 wire net1391;
 wire net1392;
 wire net1393;
 wire net1394;
 wire net1395;
 wire net1396;
 wire net1397;
 wire net1398;
 wire net1399;
 wire net14;
 wire net140;
 wire net1400;
 wire net1401;
 wire net1402;
 wire net1403;
 wire net1404;
 wire net1405;
 wire net1406;
 wire net1407;
 wire net1408;
 wire net1409;
 wire net141;
 wire net1410;
 wire net1411;
 wire net1412;
 wire net1413;
 wire net1414;
 wire net1415;
 wire net1416;
 wire net1417;
 wire net1418;
 wire net1419;
 wire net142;
 wire net1420;
 wire net1421;
 wire net1422;
 wire net1423;
 wire net1424;
 wire net1425;
 wire net1426;
 wire net1427;
 wire net1428;
 wire net1429;
 wire net143;
 wire net1430;
 wire net1431;
 wire net1432;
 wire net1433;
 wire net1434;
 wire net1435;
 wire net1436;
 wire net1437;
 wire net1438;
 wire net1439;
 wire net144;
 wire net1440;
 wire net1441;
 wire net1442;
 wire net1443;
 wire net1444;
 wire net1445;
 wire net1446;
 wire net1447;
 wire net1448;
 wire net1449;
 wire net145;
 wire net1450;
 wire net1451;
 wire net1452;
 wire net1453;
 wire net1454;
 wire net1455;
 wire net1456;
 wire net1457;
 wire net1458;
 wire net1459;
 wire net146;
 wire net1460;
 wire net1461;
 wire net1462;
 wire net1463;
 wire net1464;
 wire net1465;
 wire net1466;
 wire net1467;
 wire net1468;
 wire net1469;
 wire net147;
 wire net1470;
 wire net1471;
 wire net1472;
 wire net1473;
 wire net1474;
 wire net1475;
 wire net1476;
 wire net1477;
 wire net1478;
 wire net1479;
 wire net148;
 wire net1480;
 wire net1481;
 wire net1482;
 wire net1483;
 wire net1484;
 wire net1485;
 wire net1486;
 wire net1487;
 wire net1488;
 wire net1489;
 wire net149;
 wire net1490;
 wire net1491;
 wire net1492;
 wire net1493;
 wire net1494;
 wire net1495;
 wire net1496;
 wire net1497;
 wire net1498;
 wire net1499;
 wire net15;
 wire net150;
 wire net1500;
 wire net1501;
 wire net1502;
 wire net1503;
 wire net1504;
 wire net1505;
 wire net1506;
 wire net1507;
 wire net1508;
 wire net1509;
 wire net151;
 wire net1510;
 wire net1511;
 wire net1512;
 wire net1513;
 wire net1514;
 wire net1515;
 wire net1516;
 wire net1517;
 wire net1518;
 wire net1519;
 wire net152;
 wire net1520;
 wire net1521;
 wire net1522;
 wire net1523;
 wire net1524;
 wire net1525;
 wire net1526;
 wire net1527;
 wire net1528;
 wire net1529;
 wire net153;
 wire net1530;
 wire net1531;
 wire net1532;
 wire net1533;
 wire net1534;
 wire net1535;
 wire net1536;
 wire net1537;
 wire net1538;
 wire net1539;
 wire net154;
 wire net1540;
 wire net1541;
 wire net1542;
 wire net1543;
 wire net1544;
 wire net1545;
 wire net1546;
 wire net1547;
 wire net1548;
 wire net1549;
 wire net155;
 wire net1550;
 wire net1551;
 wire net1552;
 wire net1553;
 wire net1554;
 wire net1555;
 wire net1556;
 wire net1557;
 wire net1558;
 wire net1559;
 wire net156;
 wire net1560;
 wire net1561;
 wire net1562;
 wire net1563;
 wire net1564;
 wire net1565;
 wire net1566;
 wire net1567;
 wire net1568;
 wire net1569;
 wire net157;
 wire net1570;
 wire net1571;
 wire net1572;
 wire net1573;
 wire net1574;
 wire net1575;
 wire net1576;
 wire net1577;
 wire net1578;
 wire net1579;
 wire net158;
 wire net1580;
 wire net1581;
 wire net1582;
 wire net1583;
 wire net1584;
 wire net1585;
 wire net1586;
 wire net1587;
 wire net1588;
 wire net1589;
 wire net159;
 wire net1590;
 wire net1591;
 wire net1592;
 wire net1593;
 wire net1594;
 wire net1595;
 wire net1596;
 wire net1597;
 wire net1598;
 wire net1599;
 wire net16;
 wire net160;
 wire net1600;
 wire net1601;
 wire net1602;
 wire net1603;
 wire net1604;
 wire net1605;
 wire net1606;
 wire net1607;
 wire net1608;
 wire net1609;
 wire net161;
 wire net1610;
 wire net1611;
 wire net1612;
 wire net1613;
 wire net1614;
 wire net1615;
 wire net1616;
 wire net1617;
 wire net1618;
 wire net1619;
 wire net162;
 wire net1620;
 wire net1621;
 wire net1622;
 wire net1623;
 wire net1624;
 wire net1625;
 wire net1626;
 wire net1627;
 wire net1628;
 wire net1629;
 wire net163;
 wire net1630;
 wire net1631;
 wire net1632;
 wire net1633;
 wire net1634;
 wire net1635;
 wire net1636;
 wire net1637;
 wire net1638;
 wire net1639;
 wire net164;
 wire net1640;
 wire net1641;
 wire net1642;
 wire net1643;
 wire net1644;
 wire net1645;
 wire net1646;
 wire net1647;
 wire net1648;
 wire net1649;
 wire net165;
 wire net1650;
 wire net1651;
 wire net166;
 wire net167;
 wire net168;
 wire net169;
 wire net17;
 wire net170;
 wire net171;
 wire net172;
 wire net173;
 wire net174;
 wire net175;
 wire net176;
 wire net177;
 wire net178;
 wire net179;
 wire net18;
 wire net180;
 wire net181;
 wire net182;
 wire net183;
 wire net184;
 wire net185;
 wire net186;
 wire net187;
 wire net188;
 wire net189;
 wire net19;
 wire net190;
 wire net191;
 wire net192;
 wire net193;
 wire net194;
 wire net195;
 wire net196;
 wire net197;
 wire net198;
 wire net199;
 wire net2;
 wire net20;
 wire net200;
 wire net201;
 wire net202;
 wire net203;
 wire net204;
 wire net205;
 wire net206;
 wire net207;
 wire net208;
 wire net209;
 wire net21;
 wire net210;
 wire net211;
 wire net212;
 wire net213;
 wire net214;
 wire net215;
 wire net216;
 wire net217;
 wire net218;
 wire net219;
 wire net22;
 wire net220;
 wire net221;
 wire net222;
 wire net223;
 wire net224;
 wire net225;
 wire net226;
 wire net227;
 wire net228;
 wire net229;
 wire net23;
 wire net230;
 wire net231;
 wire net232;
 wire net233;
 wire net234;
 wire net235;
 wire net236;
 wire net237;
 wire net238;
 wire net239;
 wire net24;
 wire net240;
 wire net241;
 wire net242;
 wire net243;
 wire net244;
 wire net245;
 wire net246;
 wire net247;
 wire net248;
 wire net249;
 wire net25;
 wire net250;
 wire net251;
 wire net252;
 wire net253;
 wire net254;
 wire net255;
 wire net256;
 wire net257;
 wire net258;
 wire net259;
 wire net26;
 wire net260;
 wire net261;
 wire net262;
 wire net263;
 wire net264;
 wire net265;
 wire net266;
 wire net267;
 wire net268;
 wire net269;
 wire net27;
 wire net270;
 wire net271;
 wire net272;
 wire net273;
 wire net274;
 wire net275;
 wire net276;
 wire net277;
 wire net278;
 wire net279;
 wire net28;
 wire net280;
 wire net281;
 wire net282;
 wire net283;
 wire net284;
 wire net285;
 wire net286;
 wire net287;
 wire net288;
 wire net289;
 wire net29;
 wire net290;
 wire net291;
 wire net292;
 wire net293;
 wire net294;
 wire net295;
 wire net296;
 wire net297;
 wire net298;
 wire net299;
 wire net3;
 wire net30;
 wire net300;
 wire net301;
 wire net302;
 wire net303;
 wire net304;
 wire net305;
 wire net306;
 wire net307;
 wire net308;
 wire net309;
 wire net31;
 wire net310;
 wire net311;
 wire net312;
 wire net313;
 wire net314;
 wire net315;
 wire net316;
 wire net317;
 wire net318;
 wire net319;
 wire net32;
 wire net320;
 wire net321;
 wire net322;
 wire net323;
 wire net324;
 wire net325;
 wire net326;
 wire net327;
 wire net328;
 wire net329;
 wire net33;
 wire net330;
 wire net331;
 wire net332;
 wire net333;
 wire net334;
 wire net335;
 wire net336;
 wire net337;
 wire net338;
 wire net339;
 wire net34;
 wire net340;
 wire net341;
 wire net342;
 wire net343;
 wire net344;
 wire net345;
 wire net346;
 wire net347;
 wire net348;
 wire net349;
 wire net35;
 wire net350;
 wire net351;
 wire net352;
 wire net353;
 wire net354;
 wire net355;
 wire net356;
 wire net357;
 wire net358;
 wire net359;
 wire net36;
 wire net360;
 wire net361;
 wire net362;
 wire net363;
 wire net364;
 wire net365;
 wire net366;
 wire net367;
 wire net368;
 wire net369;
 wire net37;
 wire net370;
 wire net371;
 wire net372;
 wire net373;
 wire net374;
 wire net375;
 wire net376;
 wire net377;
 wire net378;
 wire net379;
 wire net38;
 wire net380;
 wire net381;
 wire net382;
 wire net383;
 wire net384;
 wire net385;
 wire net386;
 wire net387;
 wire net388;
 wire net389;
 wire net39;
 wire net390;
 wire net391;
 wire net392;
 wire net393;
 wire net394;
 wire net395;
 wire net396;
 wire net397;
 wire net398;
 wire net399;
 wire net4;
 wire net40;
 wire net400;
 wire net401;
 wire net402;
 wire net403;
 wire net404;
 wire net405;
 wire net406;
 wire net407;
 wire net408;
 wire net409;
 wire net41;
 wire net410;
 wire net411;
 wire net412;
 wire net413;
 wire net414;
 wire net415;
 wire net416;
 wire net417;
 wire net418;
 wire net419;
 wire net42;
 wire net420;
 wire net421;
 wire net422;
 wire net423;
 wire net424;
 wire net425;
 wire net426;
 wire net427;
 wire net428;
 wire net429;
 wire net43;
 wire net430;
 wire net431;
 wire net432;
 wire net433;
 wire net434;
 wire net435;
 wire net436;
 wire net437;
 wire net438;
 wire net439;
 wire net44;
 wire net440;
 wire net441;
 wire net442;
 wire net443;
 wire net444;
 wire net445;
 wire net446;
 wire net447;
 wire net448;
 wire net449;
 wire net45;
 wire net450;
 wire net451;
 wire net452;
 wire net453;
 wire net454;
 wire net455;
 wire net456;
 wire net457;
 wire net458;
 wire net459;
 wire net46;
 wire net460;
 wire net461;
 wire net462;
 wire net463;
 wire net464;
 wire net465;
 wire net466;
 wire net467;
 wire net468;
 wire net469;
 wire net47;
 wire net470;
 wire net471;
 wire net472;
 wire net473;
 wire net474;
 wire net475;
 wire net476;
 wire net477;
 wire net478;
 wire net479;
 wire net48;
 wire net480;
 wire net481;
 wire net482;
 wire net483;
 wire net484;
 wire net485;
 wire net486;
 wire net487;
 wire net488;
 wire net489;
 wire net49;
 wire net490;
 wire net491;
 wire net492;
 wire net493;
 wire net494;
 wire net495;
 wire net496;
 wire net497;
 wire net498;
 wire net499;
 wire net5;
 wire net50;
 wire net500;
 wire net501;
 wire net502;
 wire net503;
 wire net504;
 wire net505;
 wire net506;
 wire net507;
 wire net508;
 wire net509;
 wire net51;
 wire net510;
 wire net511;
 wire net512;
 wire net513;
 wire net514;
 wire net515;
 wire net516;
 wire net517;
 wire net518;
 wire net519;
 wire net52;
 wire net520;
 wire net521;
 wire net522;
 wire net523;
 wire net524;
 wire net525;
 wire net526;
 wire net527;
 wire net528;
 wire net529;
 wire net53;
 wire net530;
 wire net531;
 wire net532;
 wire net533;
 wire net534;
 wire net535;
 wire net536;
 wire net537;
 wire net538;
 wire net539;
 wire net54;
 wire net540;
 wire net541;
 wire net542;
 wire net543;
 wire net544;
 wire net545;
 wire net546;
 wire net547;
 wire net548;
 wire net549;
 wire net55;
 wire net550;
 wire net551;
 wire net552;
 wire net553;
 wire net554;
 wire net555;
 wire net556;
 wire net557;
 wire net558;
 wire net559;
 wire net56;
 wire net560;
 wire net561;
 wire net562;
 wire net563;
 wire net564;
 wire net565;
 wire net566;
 wire net567;
 wire net568;
 wire net569;
 wire net57;
 wire net570;
 wire net571;
 wire net572;
 wire net573;
 wire net574;
 wire net575;
 wire net576;
 wire net577;
 wire net578;
 wire net579;
 wire net58;
 wire net580;
 wire net581;
 wire net582;
 wire net583;
 wire net584;
 wire net585;
 wire net586;
 wire net587;
 wire net588;
 wire net589;
 wire net59;
 wire net590;
 wire net591;
 wire net592;
 wire net593;
 wire net594;
 wire net595;
 wire net596;
 wire net597;
 wire net598;
 wire net599;
 wire net6;
 wire net60;
 wire net600;
 wire net601;
 wire net602;
 wire net603;
 wire net604;
 wire net605;
 wire net606;
 wire net607;
 wire net608;
 wire net609;
 wire net61;
 wire net610;
 wire net611;
 wire net612;
 wire net613;
 wire net614;
 wire net615;
 wire net616;
 wire net617;
 wire net62;
 wire net63;
 wire net64;
 wire net65;
 wire net658;
 wire net659;
 wire net66;
 wire net660;
 wire net661;
 wire net662;
 wire net663;
 wire net664;
 wire net665;
 wire net666;
 wire net667;
 wire net668;
 wire net669;
 wire net67;
 wire net670;
 wire net671;
 wire net672;
 wire net673;
 wire net674;
 wire net675;
 wire net676;
 wire net677;
 wire net678;
 wire net679;
 wire net68;
 wire net680;
 wire net681;
 wire net682;
 wire net683;
 wire net684;
 wire net685;
 wire net686;
 wire net687;
 wire net688;
 wire net689;
 wire net69;
 wire net690;
 wire net691;
 wire net692;
 wire net693;
 wire net694;
 wire net695;
 wire net696;
 wire net697;
 wire net698;
 wire net699;
 wire net7;
 wire net70;
 wire net700;
 wire net701;
 wire net702;
 wire net703;
 wire net704;
 wire net705;
 wire net706;
 wire net707;
 wire net708;
 wire net709;
 wire net71;
 wire net710;
 wire net711;
 wire net712;
 wire net713;
 wire net714;
 wire net715;
 wire net716;
 wire net717;
 wire net718;
 wire net719;
 wire net72;
 wire net720;
 wire net721;
 wire net722;
 wire net723;
 wire net724;
 wire net725;
 wire net726;
 wire net727;
 wire net728;
 wire net729;
 wire net73;
 wire net730;
 wire net731;
 wire net732;
 wire net733;
 wire net734;
 wire net735;
 wire net736;
 wire net737;
 wire net738;
 wire net739;
 wire net74;
 wire net740;
 wire net741;
 wire net742;
 wire net743;
 wire net744;
 wire net745;
 wire net746;
 wire net747;
 wire net748;
 wire net749;
 wire net75;
 wire net750;
 wire net751;
 wire net752;
 wire net753;
 wire net754;
 wire net755;
 wire net756;
 wire net757;
 wire net758;
 wire net759;
 wire net76;
 wire net760;
 wire net761;
 wire net762;
 wire net763;
 wire net764;
 wire net765;
 wire net766;
 wire net767;
 wire net768;
 wire net769;
 wire net77;
 wire net770;
 wire net771;
 wire net772;
 wire net773;
 wire net774;
 wire net775;
 wire net776;
 wire net777;
 wire net778;
 wire net779;
 wire net78;
 wire net780;
 wire net781;
 wire net782;
 wire net783;
 wire net784;
 wire net785;
 wire net786;
 wire net787;
 wire net788;
 wire net789;
 wire net79;
 wire net790;
 wire net791;
 wire net792;
 wire net793;
 wire net794;
 wire net795;
 wire net796;
 wire net797;
 wire net798;
 wire net799;
 wire net8;
 wire net80;
 wire net800;
 wire net801;
 wire net802;
 wire net803;
 wire net804;
 wire net805;
 wire net806;
 wire net807;
 wire net808;
 wire net809;
 wire net81;
 wire net810;
 wire net811;
 wire net812;
 wire net813;
 wire net814;
 wire net815;
 wire net816;
 wire net817;
 wire net818;
 wire net819;
 wire net82;
 wire net820;
 wire net821;
 wire net822;
 wire net823;
 wire net824;
 wire net825;
 wire net826;
 wire net827;
 wire net828;
 wire net829;
 wire net83;
 wire net830;
 wire net831;
 wire net832;
 wire net833;
 wire net834;
 wire net835;
 wire net836;
 wire net837;
 wire net838;
 wire net839;
 wire net84;
 wire net840;
 wire net841;
 wire net842;
 wire net843;
 wire net844;
 wire net845;
 wire net846;
 wire net847;
 wire net848;
 wire net849;
 wire net85;
 wire net850;
 wire net851;
 wire net852;
 wire net853;
 wire net854;
 wire net855;
 wire net856;
 wire net857;
 wire net858;
 wire net859;
 wire net86;
 wire net860;
 wire net861;
 wire net862;
 wire net863;
 wire net864;
 wire net865;
 wire net866;
 wire net867;
 wire net868;
 wire net869;
 wire net87;
 wire net870;
 wire net871;
 wire net872;
 wire net873;
 wire net874;
 wire net875;
 wire net876;
 wire net877;
 wire net878;
 wire net879;
 wire net88;
 wire net880;
 wire net881;
 wire net882;
 wire net883;
 wire net884;
 wire net885;
 wire net886;
 wire net887;
 wire net888;
 wire net889;
 wire net89;
 wire net890;
 wire net891;
 wire net892;
 wire net893;
 wire net894;
 wire net895;
 wire net896;
 wire net897;
 wire net898;
 wire net899;
 wire net9;
 wire net90;
 wire net900;
 wire net901;
 wire net902;
 wire net903;
 wire net904;
 wire net905;
 wire net906;
 wire net907;
 wire net908;
 wire net909;
 wire net91;
 wire net910;
 wire net911;
 wire net912;
 wire net913;
 wire net914;
 wire net915;
 wire net916;
 wire net917;
 wire net918;
 wire net919;
 wire net92;
 wire net920;
 wire net921;
 wire net922;
 wire net923;
 wire net924;
 wire net925;
 wire net926;
 wire net927;
 wire net928;
 wire net929;
 wire net93;
 wire net930;
 wire net931;
 wire net932;
 wire net933;
 wire net934;
 wire net935;
 wire net936;
 wire net937;
 wire net938;
 wire net939;
 wire net94;
 wire net940;
 wire net941;
 wire net942;
 wire net943;
 wire net944;
 wire net945;
 wire net946;
 wire net947;
 wire net948;
 wire net949;
 wire net95;
 wire net950;
 wire net951;
 wire net952;
 wire net953;
 wire net954;
 wire net955;
 wire net956;
 wire net957;
 wire net958;
 wire net959;
 wire net96;
 wire net960;
 wire net961;
 wire net962;
 wire net963;
 wire net964;
 wire net965;
 wire net966;
 wire net967;
 wire net968;
 wire net969;
 wire net97;
 wire net970;
 wire net971;
 wire net972;
 wire net973;
 wire net974;
 wire net975;
 wire net976;
 wire net977;
 wire net978;
 wire net979;
 wire net98;
 wire net980;
 wire net981;
 wire net982;
 wire net983;
 wire net984;
 wire net985;
 wire net986;
 wire net987;
 wire net988;
 wire net989;
 wire net99;
 wire net990;
 wire net991;
 wire net992;
 wire net993;
 wire net994;
 wire net995;
 wire net996;
 wire net997;
 wire net998;
 wire net999;
 wire \next_state[0] ;
 wire \next_state[1] ;
 wire \reg_temp[0] ;
 wire \reg_temp[100] ;
 wire \reg_temp[101] ;
 wire \reg_temp[102] ;
 wire \reg_temp[103] ;
 wire \reg_temp[104] ;
 wire \reg_temp[105] ;
 wire \reg_temp[106] ;
 wire \reg_temp[107] ;
 wire \reg_temp[108] ;
 wire \reg_temp[109] ;
 wire \reg_temp[10] ;
 wire \reg_temp[110] ;
 wire \reg_temp[111] ;
 wire \reg_temp[112] ;
 wire \reg_temp[113] ;
 wire \reg_temp[114] ;
 wire \reg_temp[115] ;
 wire \reg_temp[116] ;
 wire \reg_temp[117] ;
 wire \reg_temp[118] ;
 wire \reg_temp[119] ;
 wire \reg_temp[11] ;
 wire \reg_temp[120] ;
 wire \reg_temp[121] ;
 wire \reg_temp[122] ;
 wire \reg_temp[123] ;
 wire \reg_temp[124] ;
 wire \reg_temp[125] ;
 wire \reg_temp[126] ;
 wire \reg_temp[127] ;
 wire \reg_temp[128] ;
 wire \reg_temp[129] ;
 wire \reg_temp[12] ;
 wire \reg_temp[130] ;
 wire \reg_temp[131] ;
 wire \reg_temp[132] ;
 wire \reg_temp[133] ;
 wire \reg_temp[134] ;
 wire \reg_temp[135] ;
 wire \reg_temp[136] ;
 wire \reg_temp[137] ;
 wire \reg_temp[138] ;
 wire \reg_temp[139] ;
 wire \reg_temp[13] ;
 wire \reg_temp[140] ;
 wire \reg_temp[141] ;
 wire \reg_temp[142] ;
 wire \reg_temp[143] ;
 wire \reg_temp[144] ;
 wire \reg_temp[145] ;
 wire \reg_temp[146] ;
 wire \reg_temp[147] ;
 wire \reg_temp[148] ;
 wire \reg_temp[149] ;
 wire \reg_temp[14] ;
 wire \reg_temp[150] ;
 wire \reg_temp[151] ;
 wire \reg_temp[152] ;
 wire \reg_temp[153] ;
 wire \reg_temp[154] ;
 wire \reg_temp[155] ;
 wire \reg_temp[156] ;
 wire \reg_temp[157] ;
 wire \reg_temp[158] ;
 wire \reg_temp[159] ;
 wire \reg_temp[15] ;
 wire \reg_temp[160] ;
 wire \reg_temp[161] ;
 wire \reg_temp[162] ;
 wire \reg_temp[16] ;
 wire \reg_temp[17] ;
 wire \reg_temp[18] ;
 wire \reg_temp[19] ;
 wire \reg_temp[1] ;
 wire \reg_temp[20] ;
 wire \reg_temp[21] ;
 wire \reg_temp[22] ;
 wire \reg_temp[23] ;
 wire \reg_temp[24] ;
 wire \reg_temp[25] ;
 wire \reg_temp[26] ;
 wire \reg_temp[27] ;
 wire \reg_temp[28] ;
 wire \reg_temp[29] ;
 wire \reg_temp[2] ;
 wire \reg_temp[30] ;
 wire \reg_temp[31] ;
 wire \reg_temp[32] ;
 wire \reg_temp[33] ;
 wire \reg_temp[34] ;
 wire \reg_temp[35] ;
 wire \reg_temp[36] ;
 wire \reg_temp[37] ;
 wire \reg_temp[38] ;
 wire \reg_temp[39] ;
 wire \reg_temp[3] ;
 wire \reg_temp[40] ;
 wire \reg_temp[41] ;
 wire \reg_temp[42] ;
 wire \reg_temp[43] ;
 wire \reg_temp[44] ;
 wire \reg_temp[45] ;
 wire \reg_temp[46] ;
 wire \reg_temp[47] ;
 wire \reg_temp[48] ;
 wire \reg_temp[49] ;
 wire \reg_temp[4] ;
 wire \reg_temp[50] ;
 wire \reg_temp[51] ;
 wire \reg_temp[52] ;
 wire \reg_temp[53] ;
 wire \reg_temp[54] ;
 wire \reg_temp[55] ;
 wire \reg_temp[56] ;
 wire \reg_temp[57] ;
 wire \reg_temp[58] ;
 wire \reg_temp[59] ;
 wire \reg_temp[5] ;
 wire \reg_temp[60] ;
 wire \reg_temp[61] ;
 wire \reg_temp[62] ;
 wire \reg_temp[63] ;
 wire \reg_temp[64] ;
 wire \reg_temp[65] ;
 wire \reg_temp[66] ;
 wire \reg_temp[67] ;
 wire \reg_temp[68] ;
 wire \reg_temp[69] ;
 wire \reg_temp[6] ;
 wire \reg_temp[70] ;
 wire \reg_temp[71] ;
 wire \reg_temp[72] ;
 wire \reg_temp[73] ;
 wire \reg_temp[74] ;
 wire \reg_temp[75] ;
 wire \reg_temp[76] ;
 wire \reg_temp[77] ;
 wire \reg_temp[78] ;
 wire \reg_temp[79] ;
 wire \reg_temp[7] ;
 wire \reg_temp[80] ;
 wire \reg_temp[81] ;
 wire \reg_temp[82] ;
 wire \reg_temp[83] ;
 wire \reg_temp[84] ;
 wire \reg_temp[85] ;
 wire \reg_temp[86] ;
 wire \reg_temp[87] ;
 wire \reg_temp[88] ;
 wire \reg_temp[89] ;
 wire \reg_temp[8] ;
 wire \reg_temp[90] ;
 wire \reg_temp[91] ;
 wire \reg_temp[92] ;
 wire \reg_temp[93] ;
 wire \reg_temp[94] ;
 wire \reg_temp[95] ;
 wire \reg_temp[96] ;
 wire \reg_temp[97] ;
 wire \reg_temp[98] ;
 wire \reg_temp[99] ;
 wire \reg_temp[9] ;
 wire updateRegs;

 sky130_fd_sc_hd__diode_2 ANTENNA_1 (.DIODE(_0814_));
 sky130_fd_sc_hd__diode_2 ANTENNA_10 (.DIODE(la_data_in[53]));
 sky130_fd_sc_hd__diode_2 ANTENNA_11 (.DIODE(net168));
 sky130_fd_sc_hd__diode_2 ANTENNA_12 (.DIODE(net191));
 sky130_fd_sc_hd__diode_2 ANTENNA_13 (.DIODE(net913));
 sky130_fd_sc_hd__diode_2 ANTENNA_14 (.DIODE(net1219));
 sky130_fd_sc_hd__diode_2 ANTENNA_15 (.DIODE(_0786_));
 sky130_fd_sc_hd__diode_2 ANTENNA_16 (.DIODE(la_data_in[30]));
 sky130_fd_sc_hd__diode_2 ANTENNA_17 (.DIODE(la_data_in[34]));
 sky130_fd_sc_hd__diode_2 ANTENNA_18 (.DIODE(la_data_in[51]));
 sky130_fd_sc_hd__diode_2 ANTENNA_19 (.DIODE(net187));
 sky130_fd_sc_hd__diode_2 ANTENNA_2 (.DIODE(la_data_in[21]));
 sky130_fd_sc_hd__diode_2 ANTENNA_20 (.DIODE(clknet_leaf_11_wb_clk_i));
 sky130_fd_sc_hd__diode_2 ANTENNA_21 (.DIODE(net699));
 sky130_fd_sc_hd__diode_2 ANTENNA_22 (.DIODE(net835));
 sky130_fd_sc_hd__diode_2 ANTENNA_23 (.DIODE(net863));
 sky130_fd_sc_hd__diode_2 ANTENNA_24 (.DIODE(la_data_in[25]));
 sky130_fd_sc_hd__diode_2 ANTENNA_25 (.DIODE(net205));
 sky130_fd_sc_hd__diode_2 ANTENNA_26 (.DIODE(net592));
 sky130_fd_sc_hd__diode_2 ANTENNA_3 (.DIODE(la_data_in[22]));
 sky130_fd_sc_hd__diode_2 ANTENNA_4 (.DIODE(la_data_in[23]));
 sky130_fd_sc_hd__diode_2 ANTENNA_5 (.DIODE(la_data_in[32]));
 sky130_fd_sc_hd__diode_2 ANTENNA_6 (.DIODE(la_data_in[40]));
 sky130_fd_sc_hd__diode_2 ANTENNA_7 (.DIODE(la_data_in[45]));
 sky130_fd_sc_hd__diode_2 ANTENNA_8 (.DIODE(la_data_in[48]));
 sky130_fd_sc_hd__diode_2 ANTENNA_9 (.DIODE(la_data_in[52]));
 sky130_fd_sc_hd__diode_2 ANTENNA__1008__B (.DIODE(_0573_));
 sky130_fd_sc_hd__diode_2 ANTENNA__1009__B1 (.DIODE(_0524_));
 sky130_fd_sc_hd__diode_2 ANTENNA__1021__A (.DIODE(net695));
 sky130_fd_sc_hd__diode_2 ANTENNA__1023__B (.DIODE(_0573_));
 sky130_fd_sc_hd__diode_2 ANTENNA__1028__S (.DIODE(net590));
 sky130_fd_sc_hd__diode_2 ANTENNA__1030__S (.DIODE(net590));
 sky130_fd_sc_hd__diode_2 ANTENNA__1032__S (.DIODE(net590));
 sky130_fd_sc_hd__diode_2 ANTENNA__1034__A1 (.DIODE(\reg_temp[77] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__1034__S (.DIODE(net590));
 sky130_fd_sc_hd__diode_2 ANTENNA__1035__B1 (.DIODE(net556));
 sky130_fd_sc_hd__diode_2 ANTENNA__1037__A2 (.DIODE(net531));
 sky130_fd_sc_hd__diode_2 ANTENNA__1037__B1 (.DIODE(net556));
 sky130_fd_sc_hd__diode_2 ANTENNA__1038__S (.DIODE(_0592_));
 sky130_fd_sc_hd__diode_2 ANTENNA__1039__B2 (.DIODE(_0599_));
 sky130_fd_sc_hd__diode_2 ANTENNA__1040__S (.DIODE(net590));
 sky130_fd_sc_hd__diode_2 ANTENNA__1042__S (.DIODE(net590));
 sky130_fd_sc_hd__diode_2 ANTENNA__1045__A2 (.DIODE(net531));
 sky130_fd_sc_hd__diode_2 ANTENNA__1045__B1 (.DIODE(net556));
 sky130_fd_sc_hd__diode_2 ANTENNA__1046__S (.DIODE(net590));
 sky130_fd_sc_hd__diode_2 ANTENNA__1048__S (.DIODE(net590));
 sky130_fd_sc_hd__diode_2 ANTENNA__1049__A2 (.DIODE(net531));
 sky130_fd_sc_hd__diode_2 ANTENNA__1049__B1 (.DIODE(net556));
 sky130_fd_sc_hd__diode_2 ANTENNA__1050__S (.DIODE(net590));
 sky130_fd_sc_hd__diode_2 ANTENNA__1052__S (.DIODE(net590));
 sky130_fd_sc_hd__diode_2 ANTENNA__1054__S (.DIODE(net590));
 sky130_fd_sc_hd__diode_2 ANTENNA__1055__A2 (.DIODE(net531));
 sky130_fd_sc_hd__diode_2 ANTENNA__1056__S (.DIODE(net590));
 sky130_fd_sc_hd__diode_2 ANTENNA__1058__S (.DIODE(net590));
 sky130_fd_sc_hd__diode_2 ANTENNA__1059__A2 (.DIODE(net533));
 sky130_fd_sc_hd__diode_2 ANTENNA__1059__B1 (.DIODE(net558));
 sky130_fd_sc_hd__diode_2 ANTENNA__1061__A2 (.DIODE(net531));
 sky130_fd_sc_hd__diode_2 ANTENNA__1061__B1 (.DIODE(net556));
 sky130_fd_sc_hd__diode_2 ANTENNA__1063__A2 (.DIODE(net533));
 sky130_fd_sc_hd__diode_2 ANTENNA__1063__B1 (.DIODE(net558));
 sky130_fd_sc_hd__diode_2 ANTENNA__1064__A0 (.DIODE(\reg_temp[144] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__1065__A2 (.DIODE(net531));
 sky130_fd_sc_hd__diode_2 ANTENNA__1065__B1 (.DIODE(net556));
 sky130_fd_sc_hd__diode_2 ANTENNA__1066__A0 (.DIODE(\reg_temp[143] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__1067__A2 (.DIODE(net531));
 sky130_fd_sc_hd__diode_2 ANTENNA__1067__B1 (.DIODE(net556));
 sky130_fd_sc_hd__diode_2 ANTENNA__1067__B2 (.DIODE(_0613_));
 sky130_fd_sc_hd__diode_2 ANTENNA__1068__A0 (.DIODE(\reg_temp[142] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__1068__A1 (.DIODE(\reg_temp[60] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__1069__A2 (.DIODE(net533));
 sky130_fd_sc_hd__diode_2 ANTENNA__1069__B1 (.DIODE(net558));
 sky130_fd_sc_hd__diode_2 ANTENNA__1070__A0 (.DIODE(\reg_temp[141] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__1071__A2 (.DIODE(net533));
 sky130_fd_sc_hd__diode_2 ANTENNA__1071__B1 (.DIODE(net558));
 sky130_fd_sc_hd__diode_2 ANTENNA__1072__A0 (.DIODE(\reg_temp[140] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__1073__A2 (.DIODE(net531));
 sky130_fd_sc_hd__diode_2 ANTENNA__1073__B1 (.DIODE(net556));
 sky130_fd_sc_hd__diode_2 ANTENNA__1074__A0 (.DIODE(\reg_temp[139] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__1074__A1 (.DIODE(\reg_temp[57] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__1075__A2 (.DIODE(net531));
 sky130_fd_sc_hd__diode_2 ANTENNA__1075__B1 (.DIODE(net556));
 sky130_fd_sc_hd__diode_2 ANTENNA__1075__B2 (.DIODE(_0617_));
 sky130_fd_sc_hd__diode_2 ANTENNA__1076__A0 (.DIODE(\reg_temp[138] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__1076__A1 (.DIODE(\reg_temp[56] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__1077__A2 (.DIODE(net531));
 sky130_fd_sc_hd__diode_2 ANTENNA__1077__B1 (.DIODE(net556));
 sky130_fd_sc_hd__diode_2 ANTENNA__1077__B2 (.DIODE(_0618_));
 sky130_fd_sc_hd__diode_2 ANTENNA__1078__A0 (.DIODE(\reg_temp[137] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__1078__A1 (.DIODE(\reg_temp[55] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__1079__A2 (.DIODE(net531));
 sky130_fd_sc_hd__diode_2 ANTENNA__1079__B1 (.DIODE(net556));
 sky130_fd_sc_hd__diode_2 ANTENNA__1079__B2 (.DIODE(_0619_));
 sky130_fd_sc_hd__diode_2 ANTENNA__1080__A0 (.DIODE(\reg_temp[136] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__1081__A2 (.DIODE(net531));
 sky130_fd_sc_hd__diode_2 ANTENNA__1081__B1 (.DIODE(net556));
 sky130_fd_sc_hd__diode_2 ANTENNA__1081__B2 (.DIODE(_0620_));
 sky130_fd_sc_hd__diode_2 ANTENNA__1082__A0 (.DIODE(\reg_temp[135] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__1082__A1 (.DIODE(\reg_temp[53] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__1083__A2 (.DIODE(net531));
 sky130_fd_sc_hd__diode_2 ANTENNA__1083__B1 (.DIODE(net556));
 sky130_fd_sc_hd__diode_2 ANTENNA__1084__A0 (.DIODE(\reg_temp[134] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__1085__A2 (.DIODE(net531));
 sky130_fd_sc_hd__diode_2 ANTENNA__1085__B1 (.DIODE(net556));
 sky130_fd_sc_hd__diode_2 ANTENNA__1086__A0 (.DIODE(\reg_temp[133] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__1086__A1 (.DIODE(\reg_temp[51] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__1087__A2 (.DIODE(net531));
 sky130_fd_sc_hd__diode_2 ANTENNA__1087__B1 (.DIODE(net556));
 sky130_fd_sc_hd__diode_2 ANTENNA__1088__A0 (.DIODE(\reg_temp[132] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__1088__A1 (.DIODE(\reg_temp[50] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__1088__S (.DIODE(net588));
 sky130_fd_sc_hd__diode_2 ANTENNA__1089__A2 (.DIODE(net533));
 sky130_fd_sc_hd__diode_2 ANTENNA__1089__B1 (.DIODE(net558));
 sky130_fd_sc_hd__diode_2 ANTENNA__1090__A1 (.DIODE(\reg_temp[49] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__1090__S (.DIODE(net590));
 sky130_fd_sc_hd__diode_2 ANTENNA__1091__A2 (.DIODE(net533));
 sky130_fd_sc_hd__diode_2 ANTENNA__1091__B1 (.DIODE(net558));
 sky130_fd_sc_hd__diode_2 ANTENNA__1092__A0 (.DIODE(\reg_temp[130] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__1092__A1 (.DIODE(\reg_temp[48] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__1092__S (.DIODE(net585));
 sky130_fd_sc_hd__diode_2 ANTENNA__1093__A2 (.DIODE(net533));
 sky130_fd_sc_hd__diode_2 ANTENNA__1093__B1 (.DIODE(net558));
 sky130_fd_sc_hd__diode_2 ANTENNA__1094__A0 (.DIODE(\reg_temp[129] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__1094__A1 (.DIODE(\reg_temp[47] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__1094__S (.DIODE(net590));
 sky130_fd_sc_hd__diode_2 ANTENNA__1095__A2 (.DIODE(net531));
 sky130_fd_sc_hd__diode_2 ANTENNA__1095__B1 (.DIODE(net556));
 sky130_fd_sc_hd__diode_2 ANTENNA__1096__A0 (.DIODE(\reg_temp[128] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__1096__S (.DIODE(net588));
 sky130_fd_sc_hd__diode_2 ANTENNA__1097__A2 (.DIODE(net533));
 sky130_fd_sc_hd__diode_2 ANTENNA__1097__B1 (.DIODE(net558));
 sky130_fd_sc_hd__diode_2 ANTENNA__1098__A0 (.DIODE(\reg_temp[127] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__1098__A1 (.DIODE(\reg_temp[45] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__1098__S (.DIODE(net588));
 sky130_fd_sc_hd__diode_2 ANTENNA__1099__A2 (.DIODE(net530));
 sky130_fd_sc_hd__diode_2 ANTENNA__1099__B1 (.DIODE(net555));
 sky130_fd_sc_hd__diode_2 ANTENNA__1100__A0 (.DIODE(\reg_temp[126] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__1100__A1 (.DIODE(\reg_temp[44] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__1100__S (.DIODE(net585));
 sky130_fd_sc_hd__diode_2 ANTENNA__1102__A0 (.DIODE(\reg_temp[125] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__1102__A1 (.DIODE(\reg_temp[43] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__1102__S (.DIODE(net588));
 sky130_fd_sc_hd__diode_2 ANTENNA__1104__A0 (.DIODE(\reg_temp[124] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__1104__A1 (.DIODE(\reg_temp[42] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__1104__S (.DIODE(net585));
 sky130_fd_sc_hd__diode_2 ANTENNA__1106__A1 (.DIODE(\reg_temp[41] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__1106__S (.DIODE(net585));
 sky130_fd_sc_hd__diode_2 ANTENNA__1108__A0 (.DIODE(\reg_temp[122] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__1108__A1 (.DIODE(\reg_temp[40] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__1108__S (.DIODE(net585));
 sky130_fd_sc_hd__diode_2 ANTENNA__1110__A0 (.DIODE(\reg_temp[121] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__1110__A1 (.DIODE(\reg_temp[39] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__1110__S (.DIODE(net588));
 sky130_fd_sc_hd__diode_2 ANTENNA__1112__A0 (.DIODE(\reg_temp[120] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__1112__A1 (.DIODE(\reg_temp[38] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__1112__S (.DIODE(net588));
 sky130_fd_sc_hd__diode_2 ANTENNA__1113__A2 (.DIODE(net529));
 sky130_fd_sc_hd__diode_2 ANTENNA__1113__B1 (.DIODE(net554));
 sky130_fd_sc_hd__diode_2 ANTENNA__1114__A0 (.DIODE(\reg_temp[119] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__1114__A1 (.DIODE(\reg_temp[37] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__1115__A1 (.DIODE(net1303));
 sky130_fd_sc_hd__diode_2 ANTENNA__1115__A2 (.DIODE(net529));
 sky130_fd_sc_hd__diode_2 ANTENNA__1115__B1 (.DIODE(net554));
 sky130_fd_sc_hd__diode_2 ANTENNA__1116__A0 (.DIODE(\reg_temp[118] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__1116__A1 (.DIODE(\reg_temp[36] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__1117__A2 (.DIODE(net529));
 sky130_fd_sc_hd__diode_2 ANTENNA__1117__B1 (.DIODE(net554));
 sky130_fd_sc_hd__diode_2 ANTENNA__1118__A0 (.DIODE(\reg_temp[117] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__1118__A1 (.DIODE(\reg_temp[35] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__1119__A2 (.DIODE(net527));
 sky130_fd_sc_hd__diode_2 ANTENNA__1119__B1 (.DIODE(net552));
 sky130_fd_sc_hd__diode_2 ANTENNA__1120__A0 (.DIODE(\reg_temp[116] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__1120__A1 (.DIODE(\reg_temp[34] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__1121__A2 (.DIODE(net527));
 sky130_fd_sc_hd__diode_2 ANTENNA__1121__B1 (.DIODE(net552));
 sky130_fd_sc_hd__diode_2 ANTENNA__1121__B2 (.DIODE(_0640_));
 sky130_fd_sc_hd__diode_2 ANTENNA__1122__A0 (.DIODE(\reg_temp[115] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__1122__A1 (.DIODE(\reg_temp[33] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__1123__A1 (.DIODE(net1304));
 sky130_fd_sc_hd__diode_2 ANTENNA__1123__A2 (.DIODE(net529));
 sky130_fd_sc_hd__diode_2 ANTENNA__1123__B1 (.DIODE(net554));
 sky130_fd_sc_hd__diode_2 ANTENNA__1124__A0 (.DIODE(\reg_temp[114] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__1124__A1 (.DIODE(\reg_temp[32] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__1125__A2 (.DIODE(net529));
 sky130_fd_sc_hd__diode_2 ANTENNA__1125__B1 (.DIODE(net554));
 sky130_fd_sc_hd__diode_2 ANTENNA__1126__A0 (.DIODE(\reg_temp[113] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__1126__A1 (.DIODE(\reg_temp[31] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__1127__A2 (.DIODE(net527));
 sky130_fd_sc_hd__diode_2 ANTENNA__1127__B1 (.DIODE(net552));
 sky130_fd_sc_hd__diode_2 ANTENNA__1127__B2 (.DIODE(_0643_));
 sky130_fd_sc_hd__diode_2 ANTENNA__1128__A0 (.DIODE(\reg_temp[112] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__1128__A1 (.DIODE(\reg_temp[30] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__1129__A2 (.DIODE(net527));
 sky130_fd_sc_hd__diode_2 ANTENNA__1129__B1 (.DIODE(net552));
 sky130_fd_sc_hd__diode_2 ANTENNA__1129__B2 (.DIODE(_0644_));
 sky130_fd_sc_hd__diode_2 ANTENNA__1130__A0 (.DIODE(\reg_temp[111] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__1130__A1 (.DIODE(\reg_temp[29] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__1132__A0 (.DIODE(\reg_temp[110] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__1132__A1 (.DIODE(\reg_temp[28] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__1133__A2 (.DIODE(net529));
 sky130_fd_sc_hd__diode_2 ANTENNA__1133__B1 (.DIODE(net555));
 sky130_fd_sc_hd__diode_2 ANTENNA__1134__A0 (.DIODE(\reg_temp[109] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__1134__A1 (.DIODE(\reg_temp[27] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__1135__A2 (.DIODE(net530));
 sky130_fd_sc_hd__diode_2 ANTENNA__1135__B1 (.DIODE(net554));
 sky130_fd_sc_hd__diode_2 ANTENNA__1136__A0 (.DIODE(\reg_temp[108] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__1136__A1 (.DIODE(\reg_temp[26] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__1138__A0 (.DIODE(\reg_temp[107] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__1138__A1 (.DIODE(\reg_temp[25] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__1140__A0 (.DIODE(\reg_temp[106] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__1140__A1 (.DIODE(\reg_temp[24] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__1141__A2 (.DIODE(net527));
 sky130_fd_sc_hd__diode_2 ANTENNA__1141__B1 (.DIODE(net552));
 sky130_fd_sc_hd__diode_2 ANTENNA__1142__A0 (.DIODE(\reg_temp[105] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__1142__A1 (.DIODE(\reg_temp[23] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__1143__A2 (.DIODE(net527));
 sky130_fd_sc_hd__diode_2 ANTENNA__1143__B1 (.DIODE(net552));
 sky130_fd_sc_hd__diode_2 ANTENNA__1144__A0 (.DIODE(\reg_temp[104] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__1144__A1 (.DIODE(\reg_temp[22] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__1145__A2 (.DIODE(net530));
 sky130_fd_sc_hd__diode_2 ANTENNA__1145__B1 (.DIODE(net555));
 sky130_fd_sc_hd__diode_2 ANTENNA__1146__A0 (.DIODE(\reg_temp[103] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__1146__A1 (.DIODE(\reg_temp[21] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__1147__A2 (.DIODE(net527));
 sky130_fd_sc_hd__diode_2 ANTENNA__1147__B1 (.DIODE(net552));
 sky130_fd_sc_hd__diode_2 ANTENNA__1147__B2 (.DIODE(_0653_));
 sky130_fd_sc_hd__diode_2 ANTENNA__1148__A0 (.DIODE(\reg_temp[102] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__1148__A1 (.DIODE(\reg_temp[20] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__1149__A2 (.DIODE(net529));
 sky130_fd_sc_hd__diode_2 ANTENNA__1149__B1 (.DIODE(net554));
 sky130_fd_sc_hd__diode_2 ANTENNA__1150__A0 (.DIODE(\reg_temp[101] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__1150__A1 (.DIODE(\reg_temp[19] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__1151__A2 (.DIODE(net529));
 sky130_fd_sc_hd__diode_2 ANTENNA__1151__B1 (.DIODE(net554));
 sky130_fd_sc_hd__diode_2 ANTENNA__1152__A0 (.DIODE(\reg_temp[100] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__1152__A1 (.DIODE(\reg_temp[18] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__1153__A1 (.DIODE(net1227));
 sky130_fd_sc_hd__diode_2 ANTENNA__1153__A2 (.DIODE(net530));
 sky130_fd_sc_hd__diode_2 ANTENNA__1153__B1 (.DIODE(net555));
 sky130_fd_sc_hd__diode_2 ANTENNA__1154__A0 (.DIODE(\reg_temp[99] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__1154__A1 (.DIODE(\reg_temp[17] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__1155__A2 (.DIODE(net527));
 sky130_fd_sc_hd__diode_2 ANTENNA__1155__B1 (.DIODE(net552));
 sky130_fd_sc_hd__diode_2 ANTENNA__1156__A0 (.DIODE(\reg_temp[98] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__1156__A1 (.DIODE(\reg_temp[16] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__1157__A2 (.DIODE(net530));
 sky130_fd_sc_hd__diode_2 ANTENNA__1157__B1 (.DIODE(net555));
 sky130_fd_sc_hd__diode_2 ANTENNA__1158__A0 (.DIODE(\reg_temp[97] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__1158__A1 (.DIODE(\reg_temp[15] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__1159__A2 (.DIODE(net527));
 sky130_fd_sc_hd__diode_2 ANTENNA__1159__B1 (.DIODE(net552));
 sky130_fd_sc_hd__diode_2 ANTENNA__1160__A0 (.DIODE(\reg_temp[96] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__1160__A1 (.DIODE(\reg_temp[14] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__1161__A2 (.DIODE(net527));
 sky130_fd_sc_hd__diode_2 ANTENNA__1161__B1 (.DIODE(net552));
 sky130_fd_sc_hd__diode_2 ANTENNA__1162__A0 (.DIODE(\reg_temp[95] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__1162__A1 (.DIODE(\reg_temp[13] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__1162__S (.DIODE(net585));
 sky130_fd_sc_hd__diode_2 ANTENNA__1163__A2 (.DIODE(net529));
 sky130_fd_sc_hd__diode_2 ANTENNA__1163__B1 (.DIODE(net554));
 sky130_fd_sc_hd__diode_2 ANTENNA__1164__A0 (.DIODE(\reg_temp[94] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__1164__A1 (.DIODE(\reg_temp[12] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__1164__S (.DIODE(net585));
 sky130_fd_sc_hd__diode_2 ANTENNA__1165__A2 (.DIODE(net529));
 sky130_fd_sc_hd__diode_2 ANTENNA__1165__B1 (.DIODE(net554));
 sky130_fd_sc_hd__diode_2 ANTENNA__1166__A1 (.DIODE(\reg_temp[11] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__1166__S (.DIODE(net585));
 sky130_fd_sc_hd__diode_2 ANTENNA__1167__A2 (.DIODE(net529));
 sky130_fd_sc_hd__diode_2 ANTENNA__1167__B1 (.DIODE(net554));
 sky130_fd_sc_hd__diode_2 ANTENNA__1168__A1 (.DIODE(\reg_temp[10] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__1168__S (.DIODE(net585));
 sky130_fd_sc_hd__diode_2 ANTENNA__1169__A2 (.DIODE(net529));
 sky130_fd_sc_hd__diode_2 ANTENNA__1169__B1 (.DIODE(net554));
 sky130_fd_sc_hd__diode_2 ANTENNA__1170__A0 (.DIODE(\reg_temp[91] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__1170__A1 (.DIODE(\reg_temp[9] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__1170__S (.DIODE(net585));
 sky130_fd_sc_hd__diode_2 ANTENNA__1171__A2 (.DIODE(net527));
 sky130_fd_sc_hd__diode_2 ANTENNA__1171__B1 (.DIODE(net552));
 sky130_fd_sc_hd__diode_2 ANTENNA__1172__A0 (.DIODE(\reg_temp[90] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__1172__A1 (.DIODE(\reg_temp[8] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__1172__S (.DIODE(net585));
 sky130_fd_sc_hd__diode_2 ANTENNA__1173__A2 (.DIODE(net529));
 sky130_fd_sc_hd__diode_2 ANTENNA__1173__B1 (.DIODE(net554));
 sky130_fd_sc_hd__diode_2 ANTENNA__1174__A0 (.DIODE(\reg_temp[89] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__1174__A1 (.DIODE(\reg_temp[7] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__1175__A2 (.DIODE(net527));
 sky130_fd_sc_hd__diode_2 ANTENNA__1175__B1 (.DIODE(net552));
 sky130_fd_sc_hd__diode_2 ANTENNA__1176__A0 (.DIODE(\reg_temp[88] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__1176__A1 (.DIODE(\reg_temp[6] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__1177__A1 (.DIODE(net1315));
 sky130_fd_sc_hd__diode_2 ANTENNA__1177__A2 (.DIODE(net529));
 sky130_fd_sc_hd__diode_2 ANTENNA__1177__B1 (.DIODE(net554));
 sky130_fd_sc_hd__diode_2 ANTENNA__1178__A0 (.DIODE(\reg_temp[87] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__1178__A1 (.DIODE(\reg_temp[5] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__1179__A2 (.DIODE(net527));
 sky130_fd_sc_hd__diode_2 ANTENNA__1179__B1 (.DIODE(net552));
 sky130_fd_sc_hd__diode_2 ANTENNA__1180__A0 (.DIODE(net1636));
 sky130_fd_sc_hd__diode_2 ANTENNA__1180__S (.DIODE(net585));
 sky130_fd_sc_hd__diode_2 ANTENNA__1181__A1 (.DIODE(net1285));
 sky130_fd_sc_hd__diode_2 ANTENNA__1181__A2 (.DIODE(net529));
 sky130_fd_sc_hd__diode_2 ANTENNA__1181__B1 (.DIODE(net554));
 sky130_fd_sc_hd__diode_2 ANTENNA__1182__A1 (.DIODE(\reg_temp[3] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__1182__S (.DIODE(net585));
 sky130_fd_sc_hd__diode_2 ANTENNA__1183__A2 (.DIODE(net529));
 sky130_fd_sc_hd__diode_2 ANTENNA__1183__B1 (.DIODE(net554));
 sky130_fd_sc_hd__diode_2 ANTENNA__1184__A0 (.DIODE(\reg_temp[84] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__1184__A1 (.DIODE(\reg_temp[2] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__1184__S (.DIODE(net585));
 sky130_fd_sc_hd__diode_2 ANTENNA__1185__A2 (.DIODE(net527));
 sky130_fd_sc_hd__diode_2 ANTENNA__1185__B1 (.DIODE(net552));
 sky130_fd_sc_hd__diode_2 ANTENNA__1186__A0 (.DIODE(\reg_temp[83] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__1186__A1 (.DIODE(\reg_temp[1] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__1186__S (.DIODE(net585));
 sky130_fd_sc_hd__diode_2 ANTENNA__1187__A2 (.DIODE(net527));
 sky130_fd_sc_hd__diode_2 ANTENNA__1187__B1 (.DIODE(net552));
 sky130_fd_sc_hd__diode_2 ANTENNA__1188__A1 (.DIODE(\reg_temp[0] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__1188__S (.DIODE(net585));
 sky130_fd_sc_hd__diode_2 ANTENNA__1189__A2 (.DIODE(net527));
 sky130_fd_sc_hd__diode_2 ANTENNA__1189__B1 (.DIODE(net552));
 sky130_fd_sc_hd__diode_2 ANTENNA__1190__A1 (.DIODE(_0524_));
 sky130_fd_sc_hd__diode_2 ANTENNA__1191__A (.DIODE(net695));
 sky130_fd_sc_hd__diode_2 ANTENNA__1193__A (.DIODE(_0524_));
 sky130_fd_sc_hd__diode_2 ANTENNA__1194__C_N (.DIODE(_0006_));
 sky130_fd_sc_hd__diode_2 ANTENNA__1195__A0 (.DIODE(net695));
 sky130_fd_sc_hd__diode_2 ANTENNA__1197__D (.DIODE(net564));
 sky130_fd_sc_hd__diode_2 ANTENNA__1202__A2 (.DIODE(net260));
 sky130_fd_sc_hd__diode_2 ANTENNA__1202__B1 (.DIODE(_0006_));
 sky130_fd_sc_hd__diode_2 ANTENNA__1204__A (.DIODE(net695));
 sky130_fd_sc_hd__diode_2 ANTENNA__1206__A1 (.DIODE(net70));
 sky130_fd_sc_hd__diode_2 ANTENNA__1206__A2 (.DIODE(net564));
 sky130_fd_sc_hd__diode_2 ANTENNA__1207__S (.DIODE(net525));
 sky130_fd_sc_hd__diode_2 ANTENNA__1209__A1 (.DIODE(net69));
 sky130_fd_sc_hd__diode_2 ANTENNA__1210__S (.DIODE(net525));
 sky130_fd_sc_hd__diode_2 ANTENNA__1212__A1 (.DIODE(net68));
 sky130_fd_sc_hd__diode_2 ANTENNA__1213__S (.DIODE(net525));
 sky130_fd_sc_hd__diode_2 ANTENNA__1215__A1 (.DIODE(net66));
 sky130_fd_sc_hd__diode_2 ANTENNA__1215__C1 (.DIODE(net955));
 sky130_fd_sc_hd__diode_2 ANTENNA__1216__S (.DIODE(net525));
 sky130_fd_sc_hd__diode_2 ANTENNA__1218__A1 (.DIODE(net65));
 sky130_fd_sc_hd__diode_2 ANTENNA__1218__A2 (.DIODE(net568));
 sky130_fd_sc_hd__diode_2 ANTENNA__1218__B1 (.DIODE(net581));
 sky130_fd_sc_hd__diode_2 ANTENNA__1218__C1 (.DIODE(net1072));
 sky130_fd_sc_hd__diode_2 ANTENNA__1219__S (.DIODE(net525));
 sky130_fd_sc_hd__diode_2 ANTENNA__1221__A1 (.DIODE(net64));
 sky130_fd_sc_hd__diode_2 ANTENNA__1221__A2 (.DIODE(net568));
 sky130_fd_sc_hd__diode_2 ANTENNA__1221__B1 (.DIODE(net581));
 sky130_fd_sc_hd__diode_2 ANTENNA__1221__C1 (.DIODE(net1172));
 sky130_fd_sc_hd__diode_2 ANTENNA__1222__S (.DIODE(net525));
 sky130_fd_sc_hd__diode_2 ANTENNA__1224__A1 (.DIODE(net63));
 sky130_fd_sc_hd__diode_2 ANTENNA__1224__A2 (.DIODE(net568));
 sky130_fd_sc_hd__diode_2 ANTENNA__1224__B1 (.DIODE(net581));
 sky130_fd_sc_hd__diode_2 ANTENNA__1224__C1 (.DIODE(net1100));
 sky130_fd_sc_hd__diode_2 ANTENNA__1225__S (.DIODE(net525));
 sky130_fd_sc_hd__diode_2 ANTENNA__1227__A1 (.DIODE(net62));
 sky130_fd_sc_hd__diode_2 ANTENNA__1227__A2 (.DIODE(net568));
 sky130_fd_sc_hd__diode_2 ANTENNA__1227__B1 (.DIODE(net581));
 sky130_fd_sc_hd__diode_2 ANTENNA__1227__C1 (.DIODE(net1079));
 sky130_fd_sc_hd__diode_2 ANTENNA__1228__S (.DIODE(net525));
 sky130_fd_sc_hd__diode_2 ANTENNA__1230__A1 (.DIODE(net61));
 sky130_fd_sc_hd__diode_2 ANTENNA__1230__A2 (.DIODE(net568));
 sky130_fd_sc_hd__diode_2 ANTENNA__1230__B1 (.DIODE(net581));
 sky130_fd_sc_hd__diode_2 ANTENNA__1230__C1 (.DIODE(net1005));
 sky130_fd_sc_hd__diode_2 ANTENNA__1231__S (.DIODE(net525));
 sky130_fd_sc_hd__diode_2 ANTENNA__1233__A1 (.DIODE(net60));
 sky130_fd_sc_hd__diode_2 ANTENNA__1233__A2 (.DIODE(net568));
 sky130_fd_sc_hd__diode_2 ANTENNA__1233__B1 (.DIODE(net581));
 sky130_fd_sc_hd__diode_2 ANTENNA__1234__S (.DIODE(net525));
 sky130_fd_sc_hd__diode_2 ANTENNA__1236__A1 (.DIODE(net59));
 sky130_fd_sc_hd__diode_2 ANTENNA__1237__S (.DIODE(net525));
 sky130_fd_sc_hd__diode_2 ANTENNA__1239__A1 (.DIODE(net58));
 sky130_fd_sc_hd__diode_2 ANTENNA__1240__S (.DIODE(net525));
 sky130_fd_sc_hd__diode_2 ANTENNA__1242__A1 (.DIODE(net57));
 sky130_fd_sc_hd__diode_2 ANTENNA__1243__S (.DIODE(net525));
 sky130_fd_sc_hd__diode_2 ANTENNA__1245__A1 (.DIODE(net55));
 sky130_fd_sc_hd__diode_2 ANTENNA__1246__S (.DIODE(net525));
 sky130_fd_sc_hd__diode_2 ANTENNA__1248__A1 (.DIODE(net54));
 sky130_fd_sc_hd__diode_2 ANTENNA__1249__S (.DIODE(net525));
 sky130_fd_sc_hd__diode_2 ANTENNA__1251__A1 (.DIODE(net53));
 sky130_fd_sc_hd__diode_2 ANTENNA__1252__S (.DIODE(net525));
 sky130_fd_sc_hd__diode_2 ANTENNA__1254__A1 (.DIODE(net52));
 sky130_fd_sc_hd__diode_2 ANTENNA__1254__A2 (.DIODE(net568));
 sky130_fd_sc_hd__diode_2 ANTENNA__1254__B1 (.DIODE(net581));
 sky130_fd_sc_hd__diode_2 ANTENNA__1255__S (.DIODE(net683));
 sky130_fd_sc_hd__diode_2 ANTENNA__1257__A1 (.DIODE(net51));
 sky130_fd_sc_hd__diode_2 ANTENNA__1257__A2 (.DIODE(net571));
 sky130_fd_sc_hd__diode_2 ANTENNA__1257__B1 (.DIODE(net584));
 sky130_fd_sc_hd__diode_2 ANTENNA__1258__S (.DIODE(net683));
 sky130_fd_sc_hd__diode_2 ANTENNA__1260__A1 (.DIODE(net50));
 sky130_fd_sc_hd__diode_2 ANTENNA__1260__A2 (.DIODE(net571));
 sky130_fd_sc_hd__diode_2 ANTENNA__1260__B1 (.DIODE(net584));
 sky130_fd_sc_hd__diode_2 ANTENNA__1261__A1 (.DIODE(\reg_temp[144] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__1261__S (.DIODE(net683));
 sky130_fd_sc_hd__diode_2 ANTENNA__1263__A1 (.DIODE(net49));
 sky130_fd_sc_hd__diode_2 ANTENNA__1263__A2 (.DIODE(net571));
 sky130_fd_sc_hd__diode_2 ANTENNA__1263__B1 (.DIODE(net584));
 sky130_fd_sc_hd__diode_2 ANTENNA__1263__B2 (.DIODE(\reg_temp[144] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__1264__S (.DIODE(net683));
 sky130_fd_sc_hd__diode_2 ANTENNA__1266__A2 (.DIODE(net571));
 sky130_fd_sc_hd__diode_2 ANTENNA__1266__B1 (.DIODE(net584));
 sky130_fd_sc_hd__diode_2 ANTENNA__1266__B2 (.DIODE(\reg_temp[143] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__1267__A1 (.DIODE(\reg_temp[142] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__1267__S (.DIODE(net683));
 sky130_fd_sc_hd__diode_2 ANTENNA__1269__A2 (.DIODE(net571));
 sky130_fd_sc_hd__diode_2 ANTENNA__1269__B1 (.DIODE(net584));
 sky130_fd_sc_hd__diode_2 ANTENNA__1269__B2 (.DIODE(\reg_temp[142] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__1270__A1 (.DIODE(\reg_temp[141] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__1270__S (.DIODE(net524));
 sky130_fd_sc_hd__diode_2 ANTENNA__1272__A2 (.DIODE(net571));
 sky130_fd_sc_hd__diode_2 ANTENNA__1272__B1 (.DIODE(net584));
 sky130_fd_sc_hd__diode_2 ANTENNA__1272__B2 (.DIODE(\reg_temp[141] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__1273__A1 (.DIODE(\reg_temp[140] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__1273__S (.DIODE(net524));
 sky130_fd_sc_hd__diode_2 ANTENNA__1275__A2 (.DIODE(net566));
 sky130_fd_sc_hd__diode_2 ANTENNA__1275__B1 (.DIODE(net579));
 sky130_fd_sc_hd__diode_2 ANTENNA__1275__B2 (.DIODE(\reg_temp[140] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__1276__S (.DIODE(net524));
 sky130_fd_sc_hd__diode_2 ANTENNA__1278__A2 (.DIODE(net571));
 sky130_fd_sc_hd__diode_2 ANTENNA__1278__B1 (.DIODE(net584));
 sky130_fd_sc_hd__diode_2 ANTENNA__1278__B2 (.DIODE(\reg_temp[139] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__1279__S (.DIODE(net524));
 sky130_fd_sc_hd__diode_2 ANTENNA__1280__A (.DIODE(net597));
 sky130_fd_sc_hd__diode_2 ANTENNA__1281__A2 (.DIODE(net567));
 sky130_fd_sc_hd__diode_2 ANTENNA__1281__B1 (.DIODE(net580));
 sky130_fd_sc_hd__diode_2 ANTENNA__1281__B2 (.DIODE(\reg_temp[138] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__1282__A1 (.DIODE(\reg_temp[137] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__1282__S (.DIODE(net683));
 sky130_fd_sc_hd__diode_2 ANTENNA__1283__A (.DIODE(net597));
 sky130_fd_sc_hd__diode_2 ANTENNA__1284__A2 (.DIODE(net566));
 sky130_fd_sc_hd__diode_2 ANTENNA__1284__B1 (.DIODE(net579));
 sky130_fd_sc_hd__diode_2 ANTENNA__1284__B2 (.DIODE(\reg_temp[137] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__1285__A1 (.DIODE(\reg_temp[136] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__1285__S (.DIODE(net524));
 sky130_fd_sc_hd__diode_2 ANTENNA__1286__A (.DIODE(net597));
 sky130_fd_sc_hd__diode_2 ANTENNA__1287__A2 (.DIODE(net566));
 sky130_fd_sc_hd__diode_2 ANTENNA__1287__B1 (.DIODE(net579));
 sky130_fd_sc_hd__diode_2 ANTENNA__1287__B2 (.DIODE(\reg_temp[136] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__1288__A1 (.DIODE(\reg_temp[135] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__1288__S (.DIODE(net524));
 sky130_fd_sc_hd__diode_2 ANTENNA__1289__A (.DIODE(net597));
 sky130_fd_sc_hd__diode_2 ANTENNA__1290__A2 (.DIODE(net566));
 sky130_fd_sc_hd__diode_2 ANTENNA__1290__B1 (.DIODE(net579));
 sky130_fd_sc_hd__diode_2 ANTENNA__1290__B2 (.DIODE(\reg_temp[135] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__1291__A1 (.DIODE(\reg_temp[134] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__1291__S (.DIODE(net524));
 sky130_fd_sc_hd__diode_2 ANTENNA__1292__A (.DIODE(net597));
 sky130_fd_sc_hd__diode_2 ANTENNA__1293__A2 (.DIODE(net566));
 sky130_fd_sc_hd__diode_2 ANTENNA__1293__B1 (.DIODE(net579));
 sky130_fd_sc_hd__diode_2 ANTENNA__1293__B2 (.DIODE(\reg_temp[134] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__1294__A1 (.DIODE(\reg_temp[133] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__1294__S (.DIODE(net524));
 sky130_fd_sc_hd__diode_2 ANTENNA__1295__A (.DIODE(net597));
 sky130_fd_sc_hd__diode_2 ANTENNA__1296__A2 (.DIODE(net566));
 sky130_fd_sc_hd__diode_2 ANTENNA__1296__B1 (.DIODE(net579));
 sky130_fd_sc_hd__diode_2 ANTENNA__1296__B2 (.DIODE(\reg_temp[133] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__1297__A1 (.DIODE(\reg_temp[132] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__1297__S (.DIODE(net524));
 sky130_fd_sc_hd__diode_2 ANTENNA__1298__A (.DIODE(net597));
 sky130_fd_sc_hd__diode_2 ANTENNA__1299__A2 (.DIODE(net566));
 sky130_fd_sc_hd__diode_2 ANTENNA__1299__B1 (.DIODE(net579));
 sky130_fd_sc_hd__diode_2 ANTENNA__1299__B2 (.DIODE(\reg_temp[132] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__1300__A1 (.DIODE(\reg_temp[131] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__1300__S (.DIODE(net524));
 sky130_fd_sc_hd__diode_2 ANTENNA__1301__A (.DIODE(net597));
 sky130_fd_sc_hd__diode_2 ANTENNA__1302__A2 (.DIODE(net564));
 sky130_fd_sc_hd__diode_2 ANTENNA__1302__B1 (.DIODE(net580));
 sky130_fd_sc_hd__diode_2 ANTENNA__1302__B2 (.DIODE(\reg_temp[131] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__1303__A1 (.DIODE(\reg_temp[130] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__1303__S (.DIODE(net524));
 sky130_fd_sc_hd__diode_2 ANTENNA__1304__A (.DIODE(net597));
 sky130_fd_sc_hd__diode_2 ANTENNA__1305__A2 (.DIODE(net567));
 sky130_fd_sc_hd__diode_2 ANTENNA__1305__B1 (.DIODE(net577));
 sky130_fd_sc_hd__diode_2 ANTENNA__1305__B2 (.DIODE(\reg_temp[130] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__1306__A1 (.DIODE(\reg_temp[129] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__1306__S (.DIODE(net524));
 sky130_fd_sc_hd__diode_2 ANTENNA__1307__A (.DIODE(net597));
 sky130_fd_sc_hd__diode_2 ANTENNA__1308__A2 (.DIODE(net564));
 sky130_fd_sc_hd__diode_2 ANTENNA__1308__B1 (.DIODE(net577));
 sky130_fd_sc_hd__diode_2 ANTENNA__1308__B2 (.DIODE(\reg_temp[129] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__1309__A1 (.DIODE(\reg_temp[128] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__1309__S (.DIODE(net524));
 sky130_fd_sc_hd__diode_2 ANTENNA__1310__A (.DIODE(net597));
 sky130_fd_sc_hd__diode_2 ANTENNA__1311__A2 (.DIODE(net564));
 sky130_fd_sc_hd__diode_2 ANTENNA__1311__B1 (.DIODE(net577));
 sky130_fd_sc_hd__diode_2 ANTENNA__1311__B2 (.DIODE(\reg_temp[128] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__1312__A1 (.DIODE(\reg_temp[127] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__1312__S (.DIODE(net524));
 sky130_fd_sc_hd__diode_2 ANTENNA__1314__A2 (.DIODE(net564));
 sky130_fd_sc_hd__diode_2 ANTENNA__1314__B1 (.DIODE(net580));
 sky130_fd_sc_hd__diode_2 ANTENNA__1314__B2 (.DIODE(\reg_temp[127] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__1315__S (.DIODE(net524));
 sky130_fd_sc_hd__diode_2 ANTENNA__1317__A2 (.DIODE(net567));
 sky130_fd_sc_hd__diode_2 ANTENNA__1317__B1 (.DIODE(net577));
 sky130_fd_sc_hd__diode_2 ANTENNA__1317__B2 (.DIODE(\reg_temp[126] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__1318__A1 (.DIODE(\reg_temp[125] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__1318__S (.DIODE(net524));
 sky130_fd_sc_hd__diode_2 ANTENNA__1320__A1 (.DIODE(net28));
 sky130_fd_sc_hd__diode_2 ANTENNA__1320__A2 (.DIODE(net567));
 sky130_fd_sc_hd__diode_2 ANTENNA__1320__B1 (.DIODE(net577));
 sky130_fd_sc_hd__diode_2 ANTENNA__1320__B2 (.DIODE(\reg_temp[125] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__1321__A1 (.DIODE(\reg_temp[124] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__1321__S (.DIODE(net684));
 sky130_fd_sc_hd__diode_2 ANTENNA__1323__A1 (.DIODE(net27));
 sky130_fd_sc_hd__diode_2 ANTENNA__1323__A2 (.DIODE(net564));
 sky130_fd_sc_hd__diode_2 ANTENNA__1323__B1 (.DIODE(net577));
 sky130_fd_sc_hd__diode_2 ANTENNA__1323__B2 (.DIODE(\reg_temp[124] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__1324__A1 (.DIODE(\reg_temp[123] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__1324__S (.DIODE(net684));
 sky130_fd_sc_hd__diode_2 ANTENNA__1326__A2 (.DIODE(net564));
 sky130_fd_sc_hd__diode_2 ANTENNA__1326__B1 (.DIODE(net577));
 sky130_fd_sc_hd__diode_2 ANTENNA__1326__B2 (.DIODE(\reg_temp[123] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__1327__A1 (.DIODE(\reg_temp[122] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__1327__S (.DIODE(net684));
 sky130_fd_sc_hd__diode_2 ANTENNA__1329__A2 (.DIODE(net564));
 sky130_fd_sc_hd__diode_2 ANTENNA__1329__B1 (.DIODE(net577));
 sky130_fd_sc_hd__diode_2 ANTENNA__1329__B2 (.DIODE(\reg_temp[122] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__1330__S (.DIODE(net684));
 sky130_fd_sc_hd__diode_2 ANTENNA__1332__A2 (.DIODE(net564));
 sky130_fd_sc_hd__diode_2 ANTENNA__1332__B1 (.DIODE(net577));
 sky130_fd_sc_hd__diode_2 ANTENNA__1332__B2 (.DIODE(\reg_temp[121] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__1333__S (.DIODE(net684));
 sky130_fd_sc_hd__diode_2 ANTENNA__1335__B2 (.DIODE(\reg_temp[120] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__1336__S (.DIODE(net684));
 sky130_fd_sc_hd__diode_2 ANTENNA__1338__B2 (.DIODE(\reg_temp[119] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__1339__A1 (.DIODE(\reg_temp[118] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__1341__B2 (.DIODE(\reg_temp[118] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__1342__A1 (.DIODE(\reg_temp[117] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__1343__A (.DIODE(net592));
 sky130_fd_sc_hd__diode_2 ANTENNA__1344__B2 (.DIODE(\reg_temp[117] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__1344__C1 (.DIODE(net793));
 sky130_fd_sc_hd__diode_2 ANTENNA__1345__S (.DIODE(net522));
 sky130_fd_sc_hd__diode_2 ANTENNA__1346__A (.DIODE(net592));
 sky130_fd_sc_hd__diode_2 ANTENNA__1347__B2 (.DIODE(\reg_temp[116] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__1347__C1 (.DIODE(net763));
 sky130_fd_sc_hd__diode_2 ANTENNA__1350__B2 (.DIODE(\reg_temp[115] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__1350__C1 (.DIODE(net1063));
 sky130_fd_sc_hd__diode_2 ANTENNA__1351__S (.DIODE(net522));
 sky130_fd_sc_hd__diode_2 ANTENNA__1352__A (.DIODE(net592));
 sky130_fd_sc_hd__diode_2 ANTENNA__1353__B1 (.DIODE(net579));
 sky130_fd_sc_hd__diode_2 ANTENNA__1353__B2 (.DIODE(\reg_temp[114] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__1353__C1 (.DIODE(net901));
 sky130_fd_sc_hd__diode_2 ANTENNA__1355__A (.DIODE(net592));
 sky130_fd_sc_hd__diode_2 ANTENNA__1356__B1 (.DIODE(net579));
 sky130_fd_sc_hd__diode_2 ANTENNA__1356__B2 (.DIODE(\reg_temp[113] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__1356__C1 (.DIODE(net933));
 sky130_fd_sc_hd__diode_2 ANTENNA__1358__A (.DIODE(net592));
 sky130_fd_sc_hd__diode_2 ANTENNA__1359__A2 (.DIODE(net566));
 sky130_fd_sc_hd__diode_2 ANTENNA__1359__B1 (.DIODE(net579));
 sky130_fd_sc_hd__diode_2 ANTENNA__1359__B2 (.DIODE(\reg_temp[112] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__1359__C1 (.DIODE(net947));
 sky130_fd_sc_hd__diode_2 ANTENNA__1360__A1 (.DIODE(\reg_temp[111] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__1361__A (.DIODE(net592));
 sky130_fd_sc_hd__diode_2 ANTENNA__1362__A2 (.DIODE(net566));
 sky130_fd_sc_hd__diode_2 ANTENNA__1362__B2 (.DIODE(\reg_temp[111] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__1362__C1 (.DIODE(net880));
 sky130_fd_sc_hd__diode_2 ANTENNA__1364__A (.DIODE(net592));
 sky130_fd_sc_hd__diode_2 ANTENNA__1365__A2 (.DIODE(net566));
 sky130_fd_sc_hd__diode_2 ANTENNA__1365__B2 (.DIODE(\reg_temp[110] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__1365__C1 (.DIODE(net894));
 sky130_fd_sc_hd__diode_2 ANTENNA__1367__A (.DIODE(net592));
 sky130_fd_sc_hd__diode_2 ANTENNA__1368__A2 (.DIODE(net566));
 sky130_fd_sc_hd__diode_2 ANTENNA__1368__B2 (.DIODE(\reg_temp[109] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__1368__C1 (.DIODE(net905));
 sky130_fd_sc_hd__diode_2 ANTENNA__1369__A1 (.DIODE(\reg_temp[108] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__1370__A (.DIODE(net592));
 sky130_fd_sc_hd__diode_2 ANTENNA__1371__B2 (.DIODE(\reg_temp[108] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__1371__C1 (.DIODE(net865));
 sky130_fd_sc_hd__diode_2 ANTENNA__1372__A1 (.DIODE(\reg_temp[107] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__1373__A (.DIODE(net592));
 sky130_fd_sc_hd__diode_2 ANTENNA__1374__B2 (.DIODE(\reg_temp[107] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__1374__C1 (.DIODE(net784));
 sky130_fd_sc_hd__diode_2 ANTENNA__1375__A1 (.DIODE(\reg_temp[106] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__1375__S (.DIODE(net522));
 sky130_fd_sc_hd__diode_2 ANTENNA__1377__B2 (.DIODE(\reg_temp[106] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__1378__S (.DIODE(net683));
 sky130_fd_sc_hd__diode_2 ANTENNA__1380__A2 (.DIODE(net566));
 sky130_fd_sc_hd__diode_2 ANTENNA__1380__B1 (.DIODE(net579));
 sky130_fd_sc_hd__diode_2 ANTENNA__1380__B2 (.DIODE(\reg_temp[105] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__1380__C1 (.DIODE(net1182));
 sky130_fd_sc_hd__diode_2 ANTENNA__1381__S (.DIODE(net522));
 sky130_fd_sc_hd__diode_2 ANTENNA__1383__B2 (.DIODE(\reg_temp[104] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__1383__C1 (.DIODE(net1186));
 sky130_fd_sc_hd__diode_2 ANTENNA__1384__S (.DIODE(net522));
 sky130_fd_sc_hd__diode_2 ANTENNA__1386__B1 (.DIODE(net579));
 sky130_fd_sc_hd__diode_2 ANTENNA__1386__B2 (.DIODE(\reg_temp[103] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__1386__C1 (.DIODE(net1178));
 sky130_fd_sc_hd__diode_2 ANTENNA__1387__S (.DIODE(net522));
 sky130_fd_sc_hd__diode_2 ANTENNA__1389__A2 (.DIODE(net563));
 sky130_fd_sc_hd__diode_2 ANTENNA__1389__B1 (.DIODE(net576));
 sky130_fd_sc_hd__diode_2 ANTENNA__1389__B2 (.DIODE(\reg_temp[102] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__1389__C1 (.DIODE(_0806_));
 sky130_fd_sc_hd__diode_2 ANTENNA__1390__S (.DIODE(net522));
 sky130_fd_sc_hd__diode_2 ANTENNA__1392__A2 (.DIODE(net563));
 sky130_fd_sc_hd__diode_2 ANTENNA__1392__B1 (.DIODE(net576));
 sky130_fd_sc_hd__diode_2 ANTENNA__1392__B2 (.DIODE(\reg_temp[101] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__1392__C1 (.DIODE(_0808_));
 sky130_fd_sc_hd__diode_2 ANTENNA__1393__S (.DIODE(net522));
 sky130_fd_sc_hd__diode_2 ANTENNA__1395__A2 (.DIODE(net563));
 sky130_fd_sc_hd__diode_2 ANTENNA__1395__B1 (.DIODE(net576));
 sky130_fd_sc_hd__diode_2 ANTENNA__1395__B2 (.DIODE(\reg_temp[100] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__1395__C1 (.DIODE(_0810_));
 sky130_fd_sc_hd__diode_2 ANTENNA__1396__S (.DIODE(net522));
 sky130_fd_sc_hd__diode_2 ANTENNA__1398__A2 (.DIODE(net566));
 sky130_fd_sc_hd__diode_2 ANTENNA__1398__B1 (.DIODE(net579));
 sky130_fd_sc_hd__diode_2 ANTENNA__1398__B2 (.DIODE(\reg_temp[99] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__1399__S (.DIODE(net522));
 sky130_fd_sc_hd__diode_2 ANTENNA__1400__A (.DIODE(net592));
 sky130_fd_sc_hd__diode_2 ANTENNA__1401__B2 (.DIODE(\reg_temp[98] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__1401__C1 (.DIODE(net789));
 sky130_fd_sc_hd__diode_2 ANTENNA__1402__S (.DIODE(net522));
 sky130_fd_sc_hd__diode_2 ANTENNA__1403__A (.DIODE(net592));
 sky130_fd_sc_hd__diode_2 ANTENNA__1404__A2 (.DIODE(net563));
 sky130_fd_sc_hd__diode_2 ANTENNA__1404__B1 (.DIODE(net576));
 sky130_fd_sc_hd__diode_2 ANTENNA__1404__B2 (.DIODE(\reg_temp[97] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__1405__S (.DIODE(net522));
 sky130_fd_sc_hd__diode_2 ANTENNA__1406__A (.DIODE(net592));
 sky130_fd_sc_hd__diode_2 ANTENNA__1407__A2 (.DIODE(_0569_));
 sky130_fd_sc_hd__diode_2 ANTENNA__1407__B1 (.DIODE(net576));
 sky130_fd_sc_hd__diode_2 ANTENNA__1407__B2 (.DIODE(\reg_temp[96] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__1408__S (.DIODE(net684));
 sky130_fd_sc_hd__diode_2 ANTENNA__1409__A (.DIODE(net592));
 sky130_fd_sc_hd__diode_2 ANTENNA__1410__A2 (.DIODE(net563));
 sky130_fd_sc_hd__diode_2 ANTENNA__1410__B1 (.DIODE(_0007_));
 sky130_fd_sc_hd__diode_2 ANTENNA__1410__B2 (.DIODE(\reg_temp[95] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__1411__A1 (.DIODE(\reg_temp[94] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__1411__S (.DIODE(net684));
 sky130_fd_sc_hd__diode_2 ANTENNA__1412__A (.DIODE(net592));
 sky130_fd_sc_hd__diode_2 ANTENNA__1413__B1 (.DIODE(net573));
 sky130_fd_sc_hd__diode_2 ANTENNA__1413__B2 (.DIODE(\reg_temp[94] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__1414__A1 (.DIODE(\reg_temp[93] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__1414__S (.DIODE(net684));
 sky130_fd_sc_hd__diode_2 ANTENNA__1415__A (.DIODE(net592));
 sky130_fd_sc_hd__diode_2 ANTENNA__1416__A2 (.DIODE(net559));
 sky130_fd_sc_hd__diode_2 ANTENNA__1416__B1 (.DIODE(net573));
 sky130_fd_sc_hd__diode_2 ANTENNA__1416__B2 (.DIODE(\reg_temp[93] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__1417__A1 (.DIODE(\reg_temp[92] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__1417__S (.DIODE(net684));
 sky130_fd_sc_hd__diode_2 ANTENNA__1419__B1 (.DIODE(net573));
 sky130_fd_sc_hd__diode_2 ANTENNA__1419__B2 (.DIODE(\reg_temp[92] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__1420__A1 (.DIODE(\reg_temp[91] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__1420__S (.DIODE(net684));
 sky130_fd_sc_hd__diode_2 ANTENNA__1422__A2 (.DIODE(net563));
 sky130_fd_sc_hd__diode_2 ANTENNA__1422__B1 (.DIODE(net576));
 sky130_fd_sc_hd__diode_2 ANTENNA__1422__B2 (.DIODE(\reg_temp[91] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__1423__A1 (.DIODE(\reg_temp[90] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__1423__S (.DIODE(net684));
 sky130_fd_sc_hd__diode_2 ANTENNA__1425__A2 (.DIODE(net563));
 sky130_fd_sc_hd__diode_2 ANTENNA__1425__B1 (.DIODE(net576));
 sky130_fd_sc_hd__diode_2 ANTENNA__1425__B2 (.DIODE(\reg_temp[90] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__1425__C1 (.DIODE(net774));
 sky130_fd_sc_hd__diode_2 ANTENNA__1426__S (.DIODE(net522));
 sky130_fd_sc_hd__diode_2 ANTENNA__1428__A2 (.DIODE(net563));
 sky130_fd_sc_hd__diode_2 ANTENNA__1428__B1 (.DIODE(net576));
 sky130_fd_sc_hd__diode_2 ANTENNA__1428__B2 (.DIODE(\reg_temp[89] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__1428__C1 (.DIODE(net721));
 sky130_fd_sc_hd__diode_2 ANTENNA__1429__A1 (.DIODE(\reg_temp[88] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__1429__S (.DIODE(net522));
 sky130_fd_sc_hd__diode_2 ANTENNA__1431__A2 (.DIODE(net563));
 sky130_fd_sc_hd__diode_2 ANTENNA__1431__B1 (.DIODE(net576));
 sky130_fd_sc_hd__diode_2 ANTENNA__1431__B2 (.DIODE(\reg_temp[88] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__1432__S (.DIODE(net522));
 sky130_fd_sc_hd__diode_2 ANTENNA__1434__A2 (.DIODE(net563));
 sky130_fd_sc_hd__diode_2 ANTENNA__1434__B1 (.DIODE(net576));
 sky130_fd_sc_hd__diode_2 ANTENNA__1434__B2 (.DIODE(\reg_temp[87] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__1435__A1 (.DIODE(net1636));
 sky130_fd_sc_hd__diode_2 ANTENNA__1435__S (.DIODE(net522));
 sky130_fd_sc_hd__diode_2 ANTENNA__1437__B1 (.DIODE(net573));
 sky130_fd_sc_hd__diode_2 ANTENNA__1437__B2 (.DIODE(\reg_temp[86] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__1438__A1 (.DIODE(\reg_temp[85] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__1438__S (.DIODE(net684));
 sky130_fd_sc_hd__diode_2 ANTENNA__1440__A2 (.DIODE(net559));
 sky130_fd_sc_hd__diode_2 ANTENNA__1440__B1 (.DIODE(net573));
 sky130_fd_sc_hd__diode_2 ANTENNA__1440__B2 (.DIODE(\reg_temp[85] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__1441__A1 (.DIODE(\reg_temp[84] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__1441__S (.DIODE(net684));
 sky130_fd_sc_hd__diode_2 ANTENNA__1443__A1 (.DIODE(net145));
 sky130_fd_sc_hd__diode_2 ANTENNA__1443__B1 (.DIODE(net573));
 sky130_fd_sc_hd__diode_2 ANTENNA__1443__B2 (.DIODE(\reg_temp[84] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__1444__A1 (.DIODE(\reg_temp[83] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__1444__S (.DIODE(net684));
 sky130_fd_sc_hd__diode_2 ANTENNA__1446__A1 (.DIODE(net144));
 sky130_fd_sc_hd__diode_2 ANTENNA__1446__B1 (.DIODE(net573));
 sky130_fd_sc_hd__diode_2 ANTENNA__1446__B2 (.DIODE(\reg_temp[83] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__1447__A1 (.DIODE(\reg_temp[82] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__1447__S (.DIODE(net684));
 sky130_fd_sc_hd__diode_2 ANTENNA__1450__B1 (.DIODE(net573));
 sky130_fd_sc_hd__diode_2 ANTENNA__1457__C1 (.DIODE(net573));
 sky130_fd_sc_hd__diode_2 ANTENNA__1459__B1 (.DIODE(_0524_));
 sky130_fd_sc_hd__diode_2 ANTENNA__1460__A1 (.DIODE(net567));
 sky130_fd_sc_hd__diode_2 ANTENNA__1460__B1 (.DIODE(net577));
 sky130_fd_sc_hd__diode_2 ANTENNA__1462__A1 (.DIODE(net567));
 sky130_fd_sc_hd__diode_2 ANTENNA__1463__A (.DIODE(\reg_temp[81] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__1465__A2 (.DIODE(net1221));
 sky130_fd_sc_hd__diode_2 ANTENNA__1466__A0 (.DIODE(_0006_));
 sky130_fd_sc_hd__diode_2 ANTENNA__1466__S (.DIODE(net1221));
 sky130_fd_sc_hd__diode_2 ANTENNA__1468__A1 (.DIODE(net597));
 sky130_fd_sc_hd__diode_2 ANTENNA__1468__B1 (.DIODE(net577));
 sky130_fd_sc_hd__diode_2 ANTENNA__1468__B2 (.DIODE(\reg_temp[82] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__1469__A1 (.DIODE(net143));
 sky130_fd_sc_hd__diode_2 ANTENNA__1469__A2 (.DIODE(net564));
 sky130_fd_sc_hd__diode_2 ANTENNA__1470__A1 (.DIODE(\reg_temp[81] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__1470__S (.DIODE(net737));
 sky130_fd_sc_hd__diode_2 ANTENNA__1471__A1 (.DIODE(net142));
 sky130_fd_sc_hd__diode_2 ANTENNA__1471__A2 (.DIODE(net564));
 sky130_fd_sc_hd__diode_2 ANTENNA__1471__B1 (.DIODE(net577));
 sky130_fd_sc_hd__diode_2 ANTENNA__1471__B2 (.DIODE(\reg_temp[81] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__1472__A0 (.DIODE(_0861_));
 sky130_fd_sc_hd__diode_2 ANTENNA__1472__S (.DIODE(net538));
 sky130_fd_sc_hd__diode_2 ANTENNA__1473__A1 (.DIODE(net140));
 sky130_fd_sc_hd__diode_2 ANTENNA__1474__S (.DIODE(net538));
 sky130_fd_sc_hd__diode_2 ANTENNA__1475__A1 (.DIODE(net139));
 sky130_fd_sc_hd__diode_2 ANTENNA__1476__S (.DIODE(net538));
 sky130_fd_sc_hd__diode_2 ANTENNA__1477__A1 (.DIODE(net138));
 sky130_fd_sc_hd__diode_2 ANTENNA__1477__C1 (.DIODE(net955));
 sky130_fd_sc_hd__diode_2 ANTENNA__1478__A1 (.DIODE(\reg_temp[77] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__1478__S (.DIODE(net538));
 sky130_fd_sc_hd__diode_2 ANTENNA__1479__A1 (.DIODE(net137));
 sky130_fd_sc_hd__diode_2 ANTENNA__1479__A2 (.DIODE(net568));
 sky130_fd_sc_hd__diode_2 ANTENNA__1479__B1 (.DIODE(net581));
 sky130_fd_sc_hd__diode_2 ANTENNA__1479__B2 (.DIODE(\reg_temp[77] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__1479__C1 (.DIODE(net1072));
 sky130_fd_sc_hd__diode_2 ANTENNA__1480__S (.DIODE(net538));
 sky130_fd_sc_hd__diode_2 ANTENNA__1481__A1 (.DIODE(net136));
 sky130_fd_sc_hd__diode_2 ANTENNA__1481__A2 (.DIODE(net568));
 sky130_fd_sc_hd__diode_2 ANTENNA__1481__B1 (.DIODE(net581));
 sky130_fd_sc_hd__diode_2 ANTENNA__1481__C1 (.DIODE(net1172));
 sky130_fd_sc_hd__diode_2 ANTENNA__1482__S (.DIODE(net538));
 sky130_fd_sc_hd__diode_2 ANTENNA__1483__A1 (.DIODE(net135));
 sky130_fd_sc_hd__diode_2 ANTENNA__1483__A2 (.DIODE(net568));
 sky130_fd_sc_hd__diode_2 ANTENNA__1483__B1 (.DIODE(net581));
 sky130_fd_sc_hd__diode_2 ANTENNA__1483__C1 (.DIODE(net1100));
 sky130_fd_sc_hd__diode_2 ANTENNA__1484__S (.DIODE(net538));
 sky130_fd_sc_hd__diode_2 ANTENNA__1485__A1 (.DIODE(net134));
 sky130_fd_sc_hd__diode_2 ANTENNA__1485__A2 (.DIODE(net568));
 sky130_fd_sc_hd__diode_2 ANTENNA__1485__B1 (.DIODE(net581));
 sky130_fd_sc_hd__diode_2 ANTENNA__1485__C1 (.DIODE(net1079));
 sky130_fd_sc_hd__diode_2 ANTENNA__1486__S (.DIODE(net538));
 sky130_fd_sc_hd__diode_2 ANTENNA__1487__A1 (.DIODE(net133));
 sky130_fd_sc_hd__diode_2 ANTENNA__1487__A2 (.DIODE(net568));
 sky130_fd_sc_hd__diode_2 ANTENNA__1487__B1 (.DIODE(net581));
 sky130_fd_sc_hd__diode_2 ANTENNA__1487__C1 (.DIODE(net1005));
 sky130_fd_sc_hd__diode_2 ANTENNA__1488__S (.DIODE(net538));
 sky130_fd_sc_hd__diode_2 ANTENNA__1489__A1 (.DIODE(net132));
 sky130_fd_sc_hd__diode_2 ANTENNA__1489__A2 (.DIODE(net568));
 sky130_fd_sc_hd__diode_2 ANTENNA__1489__B1 (.DIODE(net581));
 sky130_fd_sc_hd__diode_2 ANTENNA__1490__S (.DIODE(net538));
 sky130_fd_sc_hd__diode_2 ANTENNA__1491__A1 (.DIODE(net131));
 sky130_fd_sc_hd__diode_2 ANTENNA__1492__S (.DIODE(net539));
 sky130_fd_sc_hd__diode_2 ANTENNA__1493__A1 (.DIODE(net129));
 sky130_fd_sc_hd__diode_2 ANTENNA__1493__A2 (.DIODE(net568));
 sky130_fd_sc_hd__diode_2 ANTENNA__1493__B1 (.DIODE(net581));
 sky130_fd_sc_hd__diode_2 ANTENNA__1494__S (.DIODE(net538));
 sky130_fd_sc_hd__diode_2 ANTENNA__1495__A1 (.DIODE(net128));
 sky130_fd_sc_hd__diode_2 ANTENNA__1496__S (.DIODE(net538));
 sky130_fd_sc_hd__diode_2 ANTENNA__1497__A1 (.DIODE(net127));
 sky130_fd_sc_hd__diode_2 ANTENNA__1498__S (.DIODE(net538));
 sky130_fd_sc_hd__diode_2 ANTENNA__1499__A1 (.DIODE(net126));
 sky130_fd_sc_hd__diode_2 ANTENNA__1500__S (.DIODE(net538));
 sky130_fd_sc_hd__diode_2 ANTENNA__1501__A1 (.DIODE(net125));
 sky130_fd_sc_hd__diode_2 ANTENNA__1501__A2 (.DIODE(net568));
 sky130_fd_sc_hd__diode_2 ANTENNA__1501__B1 (.DIODE(net581));
 sky130_fd_sc_hd__diode_2 ANTENNA__1502__S (.DIODE(net538));
 sky130_fd_sc_hd__diode_2 ANTENNA__1503__A1 (.DIODE(net124));
 sky130_fd_sc_hd__diode_2 ANTENNA__1503__A2 (.DIODE(net568));
 sky130_fd_sc_hd__diode_2 ANTENNA__1503__B1 (.DIODE(net581));
 sky130_fd_sc_hd__diode_2 ANTENNA__1504__S (.DIODE(net538));
 sky130_fd_sc_hd__diode_2 ANTENNA__1505__A1 (.DIODE(net123));
 sky130_fd_sc_hd__diode_2 ANTENNA__1505__A2 (.DIODE(net571));
 sky130_fd_sc_hd__diode_2 ANTENNA__1505__B1 (.DIODE(net584));
 sky130_fd_sc_hd__diode_2 ANTENNA__1506__S (.DIODE(net539));
 sky130_fd_sc_hd__diode_2 ANTENNA__1507__A1 (.DIODE(net122));
 sky130_fd_sc_hd__diode_2 ANTENNA__1507__A2 (.DIODE(net571));
 sky130_fd_sc_hd__diode_2 ANTENNA__1507__B1 (.DIODE(net584));
 sky130_fd_sc_hd__diode_2 ANTENNA__1508__S (.DIODE(net539));
 sky130_fd_sc_hd__diode_2 ANTENNA__1509__A1 (.DIODE(net121));
 sky130_fd_sc_hd__diode_2 ANTENNA__1509__A2 (.DIODE(net571));
 sky130_fd_sc_hd__diode_2 ANTENNA__1509__B1 (.DIODE(net584));
 sky130_fd_sc_hd__diode_2 ANTENNA__1510__S (.DIODE(net539));
 sky130_fd_sc_hd__diode_2 ANTENNA__1511__A1 (.DIODE(net120));
 sky130_fd_sc_hd__diode_2 ANTENNA__1511__A2 (.DIODE(net571));
 sky130_fd_sc_hd__diode_2 ANTENNA__1511__B1 (.DIODE(net584));
 sky130_fd_sc_hd__diode_2 ANTENNA__1512__A1 (.DIODE(\reg_temp[60] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__1512__S (.DIODE(net539));
 sky130_fd_sc_hd__diode_2 ANTENNA__1513__A1 (.DIODE(net118));
 sky130_fd_sc_hd__diode_2 ANTENNA__1513__A2 (.DIODE(net571));
 sky130_fd_sc_hd__diode_2 ANTENNA__1513__B1 (.DIODE(net584));
 sky130_fd_sc_hd__diode_2 ANTENNA__1513__B2 (.DIODE(\reg_temp[60] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__1514__S (.DIODE(net539));
 sky130_fd_sc_hd__diode_2 ANTENNA__1515__A1 (.DIODE(net117));
 sky130_fd_sc_hd__diode_2 ANTENNA__1515__A2 (.DIODE(net571));
 sky130_fd_sc_hd__diode_2 ANTENNA__1515__B1 (.DIODE(net584));
 sky130_fd_sc_hd__diode_2 ANTENNA__1516__S (.DIODE(net539));
 sky130_fd_sc_hd__diode_2 ANTENNA__1517__A1 (.DIODE(net116));
 sky130_fd_sc_hd__diode_2 ANTENNA__1517__A2 (.DIODE(net566));
 sky130_fd_sc_hd__diode_2 ANTENNA__1517__B1 (.DIODE(net579));
 sky130_fd_sc_hd__diode_2 ANTENNA__1518__S (.DIODE(net539));
 sky130_fd_sc_hd__diode_2 ANTENNA__1519__A1 (.DIODE(net115));
 sky130_fd_sc_hd__diode_2 ANTENNA__1519__A2 (.DIODE(net571));
 sky130_fd_sc_hd__diode_2 ANTENNA__1519__B1 (.DIODE(net584));
 sky130_fd_sc_hd__diode_2 ANTENNA__1519__B2 (.DIODE(\reg_temp[57] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__1520__A1 (.DIODE(\reg_temp[56] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__1520__S (.DIODE(net539));
 sky130_fd_sc_hd__diode_2 ANTENNA__1521__A2 (.DIODE(net567));
 sky130_fd_sc_hd__diode_2 ANTENNA__1521__B1 (.DIODE(net580));
 sky130_fd_sc_hd__diode_2 ANTENNA__1521__B2 (.DIODE(\reg_temp[56] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__1522__A1 (.DIODE(\reg_temp[55] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__1522__S (.DIODE(net737));
 sky130_fd_sc_hd__diode_2 ANTENNA__1523__A2 (.DIODE(net567));
 sky130_fd_sc_hd__diode_2 ANTENNA__1523__B1 (.DIODE(net580));
 sky130_fd_sc_hd__diode_2 ANTENNA__1523__B2 (.DIODE(\reg_temp[55] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__1524__S (.DIODE(net737));
 sky130_fd_sc_hd__diode_2 ANTENNA__1525__A1 (.DIODE(net112));
 sky130_fd_sc_hd__diode_2 ANTENNA__1525__A2 (.DIODE(net567));
 sky130_fd_sc_hd__diode_2 ANTENNA__1525__B1 (.DIODE(net580));
 sky130_fd_sc_hd__diode_2 ANTENNA__1526__A1 (.DIODE(\reg_temp[53] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__1526__S (.DIODE(net737));
 sky130_fd_sc_hd__diode_2 ANTENNA__1527__A1 (.DIODE(net111));
 sky130_fd_sc_hd__diode_2 ANTENNA__1527__A2 (.DIODE(net567));
 sky130_fd_sc_hd__diode_2 ANTENNA__1527__B1 (.DIODE(net580));
 sky130_fd_sc_hd__diode_2 ANTENNA__1527__B2 (.DIODE(\reg_temp[53] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__1528__S (.DIODE(net737));
 sky130_fd_sc_hd__diode_2 ANTENNA__1529__A1 (.DIODE(net110));
 sky130_fd_sc_hd__diode_2 ANTENNA__1529__A2 (.DIODE(net566));
 sky130_fd_sc_hd__diode_2 ANTENNA__1529__B1 (.DIODE(net579));
 sky130_fd_sc_hd__diode_2 ANTENNA__1530__A1 (.DIODE(\reg_temp[51] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__1531__B2 (.DIODE(\reg_temp[51] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__1532__A1 (.DIODE(\reg_temp[50] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__1532__S (.DIODE(net737));
 sky130_fd_sc_hd__diode_2 ANTENNA__1533__B2 (.DIODE(\reg_temp[50] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__1534__S (.DIODE(net737));
 sky130_fd_sc_hd__diode_2 ANTENNA__1535__A1 (.DIODE(net106));
 sky130_fd_sc_hd__diode_2 ANTENNA__1535__A2 (.DIODE(net564));
 sky130_fd_sc_hd__diode_2 ANTENNA__1535__B1 (.DIODE(net577));
 sky130_fd_sc_hd__diode_2 ANTENNA__1535__B2 (.DIODE(\reg_temp[49] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__1536__A1 (.DIODE(\reg_temp[48] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__1536__S (.DIODE(net737));
 sky130_fd_sc_hd__diode_2 ANTENNA__1537__A1 (.DIODE(net105));
 sky130_fd_sc_hd__diode_2 ANTENNA__1537__A2 (.DIODE(net564));
 sky130_fd_sc_hd__diode_2 ANTENNA__1537__B1 (.DIODE(net577));
 sky130_fd_sc_hd__diode_2 ANTENNA__1537__B2 (.DIODE(\reg_temp[48] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__1538__A1 (.DIODE(\reg_temp[47] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__1538__S (.DIODE(net737));
 sky130_fd_sc_hd__diode_2 ANTENNA__1539__A1 (.DIODE(net104));
 sky130_fd_sc_hd__diode_2 ANTENNA__1539__A2 (.DIODE(net564));
 sky130_fd_sc_hd__diode_2 ANTENNA__1539__B1 (.DIODE(net577));
 sky130_fd_sc_hd__diode_2 ANTENNA__1539__B2 (.DIODE(\reg_temp[47] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__1540__A1 (.DIODE(\reg_temp[46] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__1540__S (.DIODE(net737));
 sky130_fd_sc_hd__diode_2 ANTENNA__1541__A1 (.DIODE(net103));
 sky130_fd_sc_hd__diode_2 ANTENNA__1541__A2 (.DIODE(net564));
 sky130_fd_sc_hd__diode_2 ANTENNA__1541__B1 (.DIODE(net577));
 sky130_fd_sc_hd__diode_2 ANTENNA__1541__B2 (.DIODE(\reg_temp[46] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__1542__A1 (.DIODE(\reg_temp[45] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__1542__S (.DIODE(net737));
 sky130_fd_sc_hd__diode_2 ANTENNA__1543__B1 (.DIODE(net573));
 sky130_fd_sc_hd__diode_2 ANTENNA__1543__B2 (.DIODE(\reg_temp[45] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__1544__A1 (.DIODE(\reg_temp[44] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__1544__S (.DIODE(net737));
 sky130_fd_sc_hd__diode_2 ANTENNA__1545__B1 (.DIODE(net573));
 sky130_fd_sc_hd__diode_2 ANTENNA__1545__B2 (.DIODE(\reg_temp[44] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__1547__A1 (.DIODE(net100));
 sky130_fd_sc_hd__diode_2 ANTENNA__1547__A2 (.DIODE(net559));
 sky130_fd_sc_hd__diode_2 ANTENNA__1547__B2 (.DIODE(\reg_temp[43] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__1548__A1 (.DIODE(\reg_temp[42] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__1549__A2 (.DIODE(net559));
 sky130_fd_sc_hd__diode_2 ANTENNA__1549__B2 (.DIODE(\reg_temp[42] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__1551__A2 (.DIODE(net559));
 sky130_fd_sc_hd__diode_2 ANTENNA__1551__B2 (.DIODE(\reg_temp[41] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__1553__A2 (.DIODE(net559));
 sky130_fd_sc_hd__diode_2 ANTENNA__1553__B2 (.DIODE(\reg_temp[40] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__1555__A2 (.DIODE(net559));
 sky130_fd_sc_hd__diode_2 ANTENNA__1555__B2 (.DIODE(\reg_temp[39] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__1556__S (.DIODE(net737));
 sky130_fd_sc_hd__diode_2 ANTENNA__1557__A2 (.DIODE(net561));
 sky130_fd_sc_hd__diode_2 ANTENNA__1557__B1 (.DIODE(net574));
 sky130_fd_sc_hd__diode_2 ANTENNA__1557__B2 (.DIODE(\reg_temp[38] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__1558__A1 (.DIODE(\reg_temp[37] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__1559__A2 (.DIODE(net561));
 sky130_fd_sc_hd__diode_2 ANTENNA__1559__B1 (.DIODE(net574));
 sky130_fd_sc_hd__diode_2 ANTENNA__1559__B2 (.DIODE(\reg_temp[37] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__1561__A2 (.DIODE(net561));
 sky130_fd_sc_hd__diode_2 ANTENNA__1561__B1 (.DIODE(net574));
 sky130_fd_sc_hd__diode_2 ANTENNA__1561__B2 (.DIODE(\reg_temp[36] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__1563__A2 (.DIODE(net563));
 sky130_fd_sc_hd__diode_2 ANTENNA__1563__B1 (.DIODE(net576));
 sky130_fd_sc_hd__diode_2 ANTENNA__1563__B2 (.DIODE(\reg_temp[35] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__1563__C1 (.DIODE(net793));
 sky130_fd_sc_hd__diode_2 ANTENNA__1565__A2 (.DIODE(net563));
 sky130_fd_sc_hd__diode_2 ANTENNA__1565__B1 (.DIODE(net576));
 sky130_fd_sc_hd__diode_2 ANTENNA__1565__B2 (.DIODE(\reg_temp[34] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__1565__C1 (.DIODE(net763));
 sky130_fd_sc_hd__diode_2 ANTENNA__1567__A2 (.DIODE(net563));
 sky130_fd_sc_hd__diode_2 ANTENNA__1567__B1 (.DIODE(net576));
 sky130_fd_sc_hd__diode_2 ANTENNA__1567__B2 (.DIODE(\reg_temp[33] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__1567__C1 (.DIODE(net1063));
 sky130_fd_sc_hd__diode_2 ANTENNA__1569__A2 (.DIODE(net563));
 sky130_fd_sc_hd__diode_2 ANTENNA__1569__B1 (.DIODE(net576));
 sky130_fd_sc_hd__diode_2 ANTENNA__1569__B2 (.DIODE(\reg_temp[32] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__1569__C1 (.DIODE(net901));
 sky130_fd_sc_hd__diode_2 ANTENNA__1571__A2 (.DIODE(net561));
 sky130_fd_sc_hd__diode_2 ANTENNA__1571__B1 (.DIODE(net574));
 sky130_fd_sc_hd__diode_2 ANTENNA__1571__B2 (.DIODE(\reg_temp[31] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__1571__C1 (.DIODE(net933));
 sky130_fd_sc_hd__diode_2 ANTENNA__1573__B2 (.DIODE(\reg_temp[30] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__1573__C1 (.DIODE(net947));
 sky130_fd_sc_hd__diode_2 ANTENNA__1575__B2 (.DIODE(\reg_temp[29] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__1575__C1 (.DIODE(net880));
 sky130_fd_sc_hd__diode_2 ANTENNA__1577__B2 (.DIODE(\reg_temp[28] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__1577__C1 (.DIODE(net894));
 sky130_fd_sc_hd__diode_2 ANTENNA__1579__B2 (.DIODE(\reg_temp[27] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__1579__C1 (.DIODE(net905));
 sky130_fd_sc_hd__diode_2 ANTENNA__1581__A2 (.DIODE(net561));
 sky130_fd_sc_hd__diode_2 ANTENNA__1581__B1 (.DIODE(net574));
 sky130_fd_sc_hd__diode_2 ANTENNA__1581__B2 (.DIODE(\reg_temp[26] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__1581__C1 (.DIODE(net865));
 sky130_fd_sc_hd__diode_2 ANTENNA__1583__A2 (.DIODE(net561));
 sky130_fd_sc_hd__diode_2 ANTENNA__1583__B1 (.DIODE(net574));
 sky130_fd_sc_hd__diode_2 ANTENNA__1583__B2 (.DIODE(\reg_temp[25] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__1583__C1 (.DIODE(net784));
 sky130_fd_sc_hd__diode_2 ANTENNA__1585__A2 (.DIODE(net561));
 sky130_fd_sc_hd__diode_2 ANTENNA__1585__B1 (.DIODE(net574));
 sky130_fd_sc_hd__diode_2 ANTENNA__1585__B2 (.DIODE(\reg_temp[24] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__1587__B2 (.DIODE(\reg_temp[23] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__1587__C1 (.DIODE(net1182));
 sky130_fd_sc_hd__diode_2 ANTENNA__1589__A2 (.DIODE(net561));
 sky130_fd_sc_hd__diode_2 ANTENNA__1589__B2 (.DIODE(\reg_temp[22] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__1589__C1 (.DIODE(net1186));
 sky130_fd_sc_hd__diode_2 ANTENNA__1591__A2 (.DIODE(net561));
 sky130_fd_sc_hd__diode_2 ANTENNA__1591__B1 (.DIODE(net574));
 sky130_fd_sc_hd__diode_2 ANTENNA__1591__B2 (.DIODE(\reg_temp[21] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__1591__C1 (.DIODE(net1178));
 sky130_fd_sc_hd__diode_2 ANTENNA__1593__B1 (.DIODE(net574));
 sky130_fd_sc_hd__diode_2 ANTENNA__1593__B2 (.DIODE(\reg_temp[20] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__1593__C1 (.DIODE(_0806_));
 sky130_fd_sc_hd__diode_2 ANTENNA__1595__B1 (.DIODE(net574));
 sky130_fd_sc_hd__diode_2 ANTENNA__1595__B2 (.DIODE(\reg_temp[19] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__1595__C1 (.DIODE(_0808_));
 sky130_fd_sc_hd__diode_2 ANTENNA__1597__B2 (.DIODE(\reg_temp[18] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__1597__C1 (.DIODE(_0810_));
 sky130_fd_sc_hd__diode_2 ANTENNA__1599__B2 (.DIODE(\reg_temp[17] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__1600__A1 (.DIODE(\reg_temp[16] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__1601__A2 (.DIODE(net561));
 sky130_fd_sc_hd__diode_2 ANTENNA__1601__B1 (.DIODE(net574));
 sky130_fd_sc_hd__diode_2 ANTENNA__1601__B2 (.DIODE(\reg_temp[16] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__1601__C1 (.DIODE(net789));
 sky130_fd_sc_hd__diode_2 ANTENNA__1603__A2 (.DIODE(net561));
 sky130_fd_sc_hd__diode_2 ANTENNA__1603__B1 (.DIODE(net574));
 sky130_fd_sc_hd__diode_2 ANTENNA__1603__B2 (.DIODE(\reg_temp[15] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__1604__A1 (.DIODE(\reg_temp[14] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__1605__A2 (.DIODE(net561));
 sky130_fd_sc_hd__diode_2 ANTENNA__1605__B1 (.DIODE(net574));
 sky130_fd_sc_hd__diode_2 ANTENNA__1605__B2 (.DIODE(\reg_temp[14] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__1607__A2 (.DIODE(net561));
 sky130_fd_sc_hd__diode_2 ANTENNA__1607__B1 (.DIODE(net574));
 sky130_fd_sc_hd__diode_2 ANTENNA__1607__B2 (.DIODE(\reg_temp[13] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__1609__A2 (.DIODE(net559));
 sky130_fd_sc_hd__diode_2 ANTENNA__1609__B2 (.DIODE(\reg_temp[12] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__1610__A1 (.DIODE(\reg_temp[11] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__1610__S (.DIODE(net737));
 sky130_fd_sc_hd__diode_2 ANTENNA__1611__A1 (.DIODE(net12));
 sky130_fd_sc_hd__diode_2 ANTENNA__1611__A2 (.DIODE(net559));
 sky130_fd_sc_hd__diode_2 ANTENNA__1611__B2 (.DIODE(\reg_temp[11] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__1612__A1 (.DIODE(\reg_temp[10] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__1613__A2 (.DIODE(net559));
 sky130_fd_sc_hd__diode_2 ANTENNA__1613__B2 (.DIODE(\reg_temp[10] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__1614__A1 (.DIODE(\reg_temp[9] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__1615__A2 (.DIODE(net561));
 sky130_fd_sc_hd__diode_2 ANTENNA__1615__B2 (.DIODE(\reg_temp[9] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__1617__B2 (.DIODE(\reg_temp[8] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__1617__C1 (.DIODE(net774));
 sky130_fd_sc_hd__diode_2 ANTENNA__1618__A1 (.DIODE(\reg_temp[7] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__1619__B2 (.DIODE(\reg_temp[7] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__1619__C1 (.DIODE(net721));
 sky130_fd_sc_hd__diode_2 ANTENNA__1620__A1 (.DIODE(\reg_temp[6] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__1621__A2 (.DIODE(net561));
 sky130_fd_sc_hd__diode_2 ANTENNA__1621__B1 (.DIODE(net574));
 sky130_fd_sc_hd__diode_2 ANTENNA__1621__B2 (.DIODE(\reg_temp[6] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__1623__A2 (.DIODE(net561));
 sky130_fd_sc_hd__diode_2 ANTENNA__1623__B1 (.DIODE(net574));
 sky130_fd_sc_hd__diode_2 ANTENNA__1623__B2 (.DIODE(\reg_temp[5] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__1625__A2 (.DIODE(net559));
 sky130_fd_sc_hd__diode_2 ANTENNA__1625__B2 (.DIODE(\reg_temp[4] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__1627__A2 (.DIODE(net559));
 sky130_fd_sc_hd__diode_2 ANTENNA__1627__B2 (.DIODE(\reg_temp[3] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__1628__A1 (.DIODE(\reg_temp[2] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__1629__A2 (.DIODE(net559));
 sky130_fd_sc_hd__diode_2 ANTENNA__1629__B2 (.DIODE(\reg_temp[2] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__1630__A1 (.DIODE(\reg_temp[1] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__1631__A1 (.DIODE(net1));
 sky130_fd_sc_hd__diode_2 ANTENNA__1631__A2 (.DIODE(net559));
 sky130_fd_sc_hd__diode_2 ANTENNA__1631__B2 (.DIODE(\reg_temp[1] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__1632__A1 (.DIODE(\reg_temp[0] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__1633__C (.DIODE(_0573_));
 sky130_fd_sc_hd__diode_2 ANTENNA__1637__A (.DIODE(net261));
 sky130_fd_sc_hd__diode_2 ANTENNA__1637__B (.DIODE(net559));
 sky130_fd_sc_hd__diode_2 ANTENNA__1640__B1 (.DIODE(net559));
 sky130_fd_sc_hd__diode_2 ANTENNA__1641__B (.DIODE(_0524_));
 sky130_fd_sc_hd__diode_2 ANTENNA__1642__A (.DIODE(\reg_temp[0] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__1642__B (.DIODE(net540));
 sky130_fd_sc_hd__diode_2 ANTENNA__1643__A (.DIODE(\reg_temp[1] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__1643__B (.DIODE(net540));
 sky130_fd_sc_hd__diode_2 ANTENNA__1644__A (.DIODE(\reg_temp[2] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__1644__B (.DIODE(net540));
 sky130_fd_sc_hd__diode_2 ANTENNA__1645__A (.DIODE(\reg_temp[3] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__1645__B (.DIODE(net540));
 sky130_fd_sc_hd__diode_2 ANTENNA__1646__A (.DIODE(\reg_temp[4] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__1646__B (.DIODE(net540));
 sky130_fd_sc_hd__diode_2 ANTENNA__1647__A (.DIODE(\reg_temp[5] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__1648__A (.DIODE(\reg_temp[6] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__1649__A (.DIODE(\reg_temp[7] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__1650__A (.DIODE(\reg_temp[8] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__1651__A (.DIODE(\reg_temp[9] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__1651__B (.DIODE(net540));
 sky130_fd_sc_hd__diode_2 ANTENNA__1652__A (.DIODE(\reg_temp[10] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__1652__B (.DIODE(net540));
 sky130_fd_sc_hd__diode_2 ANTENNA__1653__A (.DIODE(\reg_temp[11] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__1653__B (.DIODE(net540));
 sky130_fd_sc_hd__diode_2 ANTENNA__1654__A (.DIODE(\reg_temp[12] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__1654__B (.DIODE(net540));
 sky130_fd_sc_hd__diode_2 ANTENNA__1655__A (.DIODE(\reg_temp[13] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__1655__B (.DIODE(net540));
 sky130_fd_sc_hd__diode_2 ANTENNA__1656__A (.DIODE(\reg_temp[14] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__1657__A (.DIODE(\reg_temp[15] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__1658__A (.DIODE(\reg_temp[16] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__1659__A (.DIODE(\reg_temp[17] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__1660__A (.DIODE(\reg_temp[18] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__1661__A (.DIODE(\reg_temp[19] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__1662__A (.DIODE(\reg_temp[20] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__1663__A (.DIODE(\reg_temp[21] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__1664__A (.DIODE(\reg_temp[22] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__1665__A (.DIODE(\reg_temp[23] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__1666__A (.DIODE(\reg_temp[24] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__1667__A (.DIODE(\reg_temp[25] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__1668__A (.DIODE(\reg_temp[26] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__1669__A (.DIODE(\reg_temp[27] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__1670__A (.DIODE(\reg_temp[28] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__1671__A (.DIODE(\reg_temp[29] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__1672__A (.DIODE(\reg_temp[30] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__1673__A (.DIODE(\reg_temp[31] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__1674__A (.DIODE(\reg_temp[32] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__1675__A (.DIODE(\reg_temp[33] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__1676__A (.DIODE(\reg_temp[34] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__1677__A (.DIODE(\reg_temp[35] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__1678__A (.DIODE(\reg_temp[36] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__1679__A (.DIODE(\reg_temp[37] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__1680__A (.DIODE(\reg_temp[38] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__1681__A (.DIODE(\reg_temp[39] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__1681__B (.DIODE(net540));
 sky130_fd_sc_hd__diode_2 ANTENNA__1682__A (.DIODE(\reg_temp[40] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__1682__B (.DIODE(net543));
 sky130_fd_sc_hd__diode_2 ANTENNA__1683__A (.DIODE(\reg_temp[41] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__1683__B (.DIODE(net540));
 sky130_fd_sc_hd__diode_2 ANTENNA__1684__A (.DIODE(\reg_temp[42] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__1684__B (.DIODE(net540));
 sky130_fd_sc_hd__diode_2 ANTENNA__1685__A (.DIODE(\reg_temp[43] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__1685__B (.DIODE(net540));
 sky130_fd_sc_hd__diode_2 ANTENNA__1686__A (.DIODE(\reg_temp[44] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__1686__B (.DIODE(net540));
 sky130_fd_sc_hd__diode_2 ANTENNA__1687__A (.DIODE(\reg_temp[45] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__1687__B (.DIODE(net544));
 sky130_fd_sc_hd__diode_2 ANTENNA__1688__A (.DIODE(\reg_temp[46] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__1688__B (.DIODE(net544));
 sky130_fd_sc_hd__diode_2 ANTENNA__1689__A (.DIODE(\reg_temp[47] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__1689__B (.DIODE(net544));
 sky130_fd_sc_hd__diode_2 ANTENNA__1690__A (.DIODE(\reg_temp[48] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__1690__B (.DIODE(net544));
 sky130_fd_sc_hd__diode_2 ANTENNA__1691__A (.DIODE(\reg_temp[49] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__1691__B (.DIODE(net544));
 sky130_fd_sc_hd__diode_2 ANTENNA__1692__A (.DIODE(\reg_temp[50] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__1692__B (.DIODE(net543));
 sky130_fd_sc_hd__diode_2 ANTENNA__1693__A (.DIODE(\reg_temp[51] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__1693__B (.DIODE(net543));
 sky130_fd_sc_hd__diode_2 ANTENNA__1694__B (.DIODE(net543));
 sky130_fd_sc_hd__diode_2 ANTENNA__1695__A (.DIODE(\reg_temp[53] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__1695__B (.DIODE(net543));
 sky130_fd_sc_hd__diode_2 ANTENNA__1696__B (.DIODE(net543));
 sky130_fd_sc_hd__diode_2 ANTENNA__1697__A (.DIODE(\reg_temp[55] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__1697__B (.DIODE(net543));
 sky130_fd_sc_hd__diode_2 ANTENNA__1698__A (.DIODE(\reg_temp[56] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__1698__B (.DIODE(net543));
 sky130_fd_sc_hd__diode_2 ANTENNA__1699__A (.DIODE(\reg_temp[57] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__1699__B (.DIODE(net543));
 sky130_fd_sc_hd__diode_2 ANTENNA__1700__B (.DIODE(net543));
 sky130_fd_sc_hd__diode_2 ANTENNA__1701__B (.DIODE(net543));
 sky130_fd_sc_hd__diode_2 ANTENNA__1702__A (.DIODE(\reg_temp[60] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__1702__B (.DIODE(net543));
 sky130_fd_sc_hd__diode_2 ANTENNA__1703__B (.DIODE(net543));
 sky130_fd_sc_hd__diode_2 ANTENNA__1704__B (.DIODE(net543));
 sky130_fd_sc_hd__diode_2 ANTENNA__1705__B (.DIODE(net544));
 sky130_fd_sc_hd__diode_2 ANTENNA__1706__B (.DIODE(net543));
 sky130_fd_sc_hd__diode_2 ANTENNA__1707__B (.DIODE(net548));
 sky130_fd_sc_hd__diode_2 ANTENNA__1715__B (.DIODE(net543));
 sky130_fd_sc_hd__diode_2 ANTENNA__1718__B (.DIODE(net548));
 sky130_fd_sc_hd__diode_2 ANTENNA__1719__A (.DIODE(\reg_temp[77] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__1723__A (.DIODE(\reg_temp[81] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__1724__A (.DIODE(\reg_temp[82] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__1724__B (.DIODE(net544));
 sky130_fd_sc_hd__diode_2 ANTENNA__1725__A (.DIODE(\reg_temp[83] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__1725__B (.DIODE(net540));
 sky130_fd_sc_hd__diode_2 ANTENNA__1726__A (.DIODE(\reg_temp[84] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__1727__A (.DIODE(\reg_temp[85] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__1728__A (.DIODE(\reg_temp[86] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__1728__B (.DIODE(net548));
 sky130_fd_sc_hd__diode_2 ANTENNA__1729__A (.DIODE(\reg_temp[87] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__1729__B (.DIODE(net548));
 sky130_fd_sc_hd__diode_2 ANTENNA__1730__A (.DIODE(\reg_temp[88] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__1730__B (.DIODE(net548));
 sky130_fd_sc_hd__diode_2 ANTENNA__1731__A (.DIODE(\reg_temp[89] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__1732__A (.DIODE(\reg_temp[90] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__1733__A (.DIODE(\reg_temp[91] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__1734__A (.DIODE(\reg_temp[92] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__1735__A (.DIODE(\reg_temp[93] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__1736__A (.DIODE(\reg_temp[94] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__1737__A (.DIODE(\reg_temp[95] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__1738__A (.DIODE(\reg_temp[96] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__1738__B (.DIODE(net548));
 sky130_fd_sc_hd__diode_2 ANTENNA__1739__A (.DIODE(\reg_temp[97] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__1739__B (.DIODE(net548));
 sky130_fd_sc_hd__diode_2 ANTENNA__1740__A (.DIODE(\reg_temp[98] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__1740__B (.DIODE(net548));
 sky130_fd_sc_hd__diode_2 ANTENNA__1741__A (.DIODE(\reg_temp[99] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__1742__A (.DIODE(\reg_temp[100] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__1743__A (.DIODE(\reg_temp[101] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__1744__A (.DIODE(\reg_temp[102] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__1745__A (.DIODE(\reg_temp[103] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__1746__A (.DIODE(\reg_temp[104] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__1747__A (.DIODE(\reg_temp[105] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__1748__A (.DIODE(\reg_temp[106] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__1748__B (.DIODE(net548));
 sky130_fd_sc_hd__diode_2 ANTENNA__1749__A (.DIODE(\reg_temp[107] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__1749__B (.DIODE(net548));
 sky130_fd_sc_hd__diode_2 ANTENNA__1750__A (.DIODE(\reg_temp[108] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__1750__B (.DIODE(net548));
 sky130_fd_sc_hd__diode_2 ANTENNA__1751__A (.DIODE(\reg_temp[109] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__1751__B (.DIODE(net551));
 sky130_fd_sc_hd__diode_2 ANTENNA__1752__A (.DIODE(\reg_temp[110] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__1752__B (.DIODE(net548));
 sky130_fd_sc_hd__diode_2 ANTENNA__1753__A (.DIODE(\reg_temp[111] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__1754__A (.DIODE(\reg_temp[112] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__1755__A (.DIODE(\reg_temp[113] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__1756__A (.DIODE(\reg_temp[114] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__1757__A (.DIODE(\reg_temp[115] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__1757__B (.DIODE(net551));
 sky130_fd_sc_hd__diode_2 ANTENNA__1758__A (.DIODE(\reg_temp[116] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__1758__B (.DIODE(net548));
 sky130_fd_sc_hd__diode_2 ANTENNA__1759__A (.DIODE(\reg_temp[117] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__1759__B (.DIODE(net551));
 sky130_fd_sc_hd__diode_2 ANTENNA__1760__A (.DIODE(\reg_temp[118] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__1760__B (.DIODE(net548));
 sky130_fd_sc_hd__diode_2 ANTENNA__1761__A (.DIODE(\reg_temp[119] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__1761__B (.DIODE(net548));
 sky130_fd_sc_hd__diode_2 ANTENNA__1762__A (.DIODE(\reg_temp[120] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__1763__A (.DIODE(\reg_temp[121] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__1764__A (.DIODE(\reg_temp[122] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__1765__A (.DIODE(\reg_temp[123] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__1766__A (.DIODE(\reg_temp[124] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__1767__A (.DIODE(\reg_temp[125] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__1768__A (.DIODE(\reg_temp[126] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__1769__A (.DIODE(\reg_temp[127] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__1770__A (.DIODE(\reg_temp[128] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__1771__A (.DIODE(\reg_temp[129] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__1772__A (.DIODE(\reg_temp[130] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__1772__B (.DIODE(net551));
 sky130_fd_sc_hd__diode_2 ANTENNA__1773__A (.DIODE(\reg_temp[131] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__1774__A (.DIODE(\reg_temp[132] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__1775__A (.DIODE(\reg_temp[133] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__1776__A (.DIODE(\reg_temp[134] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__1777__A (.DIODE(\reg_temp[135] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__1778__A (.DIODE(\reg_temp[136] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__1779__A (.DIODE(\reg_temp[137] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__1780__A (.DIODE(\reg_temp[138] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__1781__A (.DIODE(\reg_temp[139] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__1782__A (.DIODE(\reg_temp[140] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__1783__A (.DIODE(\reg_temp[141] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__1784__A (.DIODE(\reg_temp[142] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__1785__A (.DIODE(\reg_temp[143] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__1786__A (.DIODE(\reg_temp[144] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__1792__B (.DIODE(net551));
 sky130_fd_sc_hd__diode_2 ANTENNA__1810__C (.DIODE(_0524_));
 sky130_fd_sc_hd__diode_2 ANTENNA__1811__A (.DIODE(_0573_));
 sky130_fd_sc_hd__diode_2 ANTENNA__1812__A (.DIODE(\reg_temp[0] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__1832__A (.DIODE(net602));
 sky130_fd_sc_hd__diode_2 ANTENNA__1833__A (.DIODE(net602));
 sky130_fd_sc_hd__diode_2 ANTENNA__1834__A (.DIODE(net602));
 sky130_fd_sc_hd__diode_2 ANTENNA__1835__A (.DIODE(net602));
 sky130_fd_sc_hd__diode_2 ANTENNA__1839__A (.DIODE(net602));
 sky130_fd_sc_hd__diode_2 ANTENNA__1840__A (.DIODE(net602));
 sky130_fd_sc_hd__diode_2 ANTENNA__1841__A (.DIODE(net602));
 sky130_fd_sc_hd__diode_2 ANTENNA__1856__A (.DIODE(net599));
 sky130_fd_sc_hd__diode_2 ANTENNA__1857__A (.DIODE(net599));
 sky130_fd_sc_hd__diode_2 ANTENNA__1858__A (.DIODE(net606));
 sky130_fd_sc_hd__diode_2 ANTENNA__1859__A (.DIODE(net606));
 sky130_fd_sc_hd__diode_2 ANTENNA__1860__A (.DIODE(net606));
 sky130_fd_sc_hd__diode_2 ANTENNA__1861__A (.DIODE(net603));
 sky130_fd_sc_hd__diode_2 ANTENNA__1862__A (.DIODE(net603));
 sky130_fd_sc_hd__diode_2 ANTENNA__1863__A (.DIODE(net603));
 sky130_fd_sc_hd__diode_2 ANTENNA__1869__A (.DIODE(net610));
 sky130_fd_sc_hd__diode_2 ANTENNA__1870__A (.DIODE(net610));
 sky130_fd_sc_hd__diode_2 ANTENNA__1871__A (.DIODE(net610));
 sky130_fd_sc_hd__diode_2 ANTENNA__1872__A (.DIODE(net610));
 sky130_fd_sc_hd__diode_2 ANTENNA__1873__A (.DIODE(net610));
 sky130_fd_sc_hd__diode_2 ANTENNA__1874__A (.DIODE(net610));
 sky130_fd_sc_hd__diode_2 ANTENNA__1875__A (.DIODE(net610));
 sky130_fd_sc_hd__diode_2 ANTENNA__1876__A (.DIODE(net610));
 sky130_fd_sc_hd__diode_2 ANTENNA__1877__A (.DIODE(net617));
 sky130_fd_sc_hd__diode_2 ANTENNA__1878__A (.DIODE(net617));
 sky130_fd_sc_hd__diode_2 ANTENNA__1879__A (.DIODE(net612));
 sky130_fd_sc_hd__diode_2 ANTENNA__1880__A (.DIODE(net613));
 sky130_fd_sc_hd__diode_2 ANTENNA__1881__A (.DIODE(net616));
 sky130_fd_sc_hd__diode_2 ANTENNA__1882__A (.DIODE(net616));
 sky130_fd_sc_hd__diode_2 ANTENNA__1883__A (.DIODE(net616));
 sky130_fd_sc_hd__diode_2 ANTENNA__1884__A (.DIODE(net617));
 sky130_fd_sc_hd__diode_2 ANTENNA__1885__A (.DIODE(net617));
 sky130_fd_sc_hd__diode_2 ANTENNA__1886__A (.DIODE(net616));
 sky130_fd_sc_hd__diode_2 ANTENNA__1887__A (.DIODE(net616));
 sky130_fd_sc_hd__diode_2 ANTENNA__1888__A (.DIODE(net617));
 sky130_fd_sc_hd__diode_2 ANTENNA__1889__A (.DIODE(net617));
 sky130_fd_sc_hd__diode_2 ANTENNA__1890__A (.DIODE(net616));
 sky130_fd_sc_hd__diode_2 ANTENNA__1894__A (.DIODE(net606));
 sky130_fd_sc_hd__diode_2 ANTENNA__1895__A (.DIODE(net613));
 sky130_fd_sc_hd__diode_2 ANTENNA__1896__A (.DIODE(net613));
 sky130_fd_sc_hd__diode_2 ANTENNA__1897__A (.DIODE(net612));
 sky130_fd_sc_hd__diode_2 ANTENNA__1898__A (.DIODE(net606));
 sky130_fd_sc_hd__diode_2 ANTENNA__1899__A (.DIODE(net606));
 sky130_fd_sc_hd__diode_2 ANTENNA__1900__A (.DIODE(net599));
 sky130_fd_sc_hd__diode_2 ANTENNA__1901__A (.DIODE(net606));
 sky130_fd_sc_hd__diode_2 ANTENNA__1902__A (.DIODE(net599));
 sky130_fd_sc_hd__diode_2 ANTENNA__1903__A (.DIODE(net599));
 sky130_fd_sc_hd__diode_2 ANTENNA__1904__A (.DIODE(net599));
 sky130_fd_sc_hd__diode_2 ANTENNA__1905__A (.DIODE(net599));
 sky130_fd_sc_hd__diode_2 ANTENNA__1908__A (.DIODE(net602));
 sky130_fd_sc_hd__diode_2 ANTENNA__1909__A (.DIODE(net602));
 sky130_fd_sc_hd__diode_2 ANTENNA__1911__A (.DIODE(net599));
 sky130_fd_sc_hd__diode_2 ANTENNA__1912__A (.DIODE(net599));
 sky130_fd_sc_hd__diode_2 ANTENNA__1913__A (.DIODE(net599));
 sky130_fd_sc_hd__diode_2 ANTENNA__1917__A (.DIODE(net603));
 sky130_fd_sc_hd__diode_2 ANTENNA__1918__A (.DIODE(net603));
 sky130_fd_sc_hd__diode_2 ANTENNA__1919__A (.DIODE(net603));
 sky130_fd_sc_hd__diode_2 ANTENNA__1920__A (.DIODE(net602));
 sky130_fd_sc_hd__diode_2 ANTENNA__1921__A (.DIODE(net602));
 sky130_fd_sc_hd__diode_2 ANTENNA__1922__A (.DIODE(net602));
 sky130_fd_sc_hd__diode_2 ANTENNA__1923__A (.DIODE(net603));
 sky130_fd_sc_hd__diode_2 ANTENNA__1924__A (.DIODE(net603));
 sky130_fd_sc_hd__diode_2 ANTENNA__1925__A (.DIODE(net603));
 sky130_fd_sc_hd__diode_2 ANTENNA__1926__A (.DIODE(net603));
 sky130_fd_sc_hd__diode_2 ANTENNA__1927__A (.DIODE(net603));
 sky130_fd_sc_hd__diode_2 ANTENNA__1928__A (.DIODE(net603));
 sky130_fd_sc_hd__diode_2 ANTENNA__1929__A (.DIODE(net603));
 sky130_fd_sc_hd__diode_2 ANTENNA__1930__A (.DIODE(net603));
 sky130_fd_sc_hd__diode_2 ANTENNA__1931__A (.DIODE(net605));
 sky130_fd_sc_hd__diode_2 ANTENNA__1936__A (.DIODE(net605));
 sky130_fd_sc_hd__diode_2 ANTENNA__1937__A (.DIODE(net605));
 sky130_fd_sc_hd__diode_2 ANTENNA__1940__A (.DIODE(net603));
 sky130_fd_sc_hd__diode_2 ANTENNA__1941__A (.DIODE(net603));
 sky130_fd_sc_hd__diode_2 ANTENNA__1942__A (.DIODE(net606));
 sky130_fd_sc_hd__diode_2 ANTENNA__1943__A (.DIODE(net606));
 sky130_fd_sc_hd__diode_2 ANTENNA__1944__A (.DIODE(net606));
 sky130_fd_sc_hd__diode_2 ANTENNA__1945__A (.DIODE(net606));
 sky130_fd_sc_hd__diode_2 ANTENNA__1946__A (.DIODE(net606));
 sky130_fd_sc_hd__diode_2 ANTENNA__1947__A (.DIODE(net606));
 sky130_fd_sc_hd__diode_2 ANTENNA__1948__A (.DIODE(net606));
 sky130_fd_sc_hd__diode_2 ANTENNA__1949__A (.DIODE(net606));
 sky130_fd_sc_hd__diode_2 ANTENNA__1955__A (.DIODE(net605));
 sky130_fd_sc_hd__diode_2 ANTENNA__1956__A (.DIODE(net605));
 sky130_fd_sc_hd__diode_2 ANTENNA__1957__A (.DIODE(net605));
 sky130_fd_sc_hd__diode_2 ANTENNA__1958__A (.DIODE(net610));
 sky130_fd_sc_hd__diode_2 ANTENNA__1959__A (.DIODE(net610));
 sky130_fd_sc_hd__diode_2 ANTENNA__1960__A (.DIODE(net610));
 sky130_fd_sc_hd__diode_2 ANTENNA__1961__A (.DIODE(net610));
 sky130_fd_sc_hd__diode_2 ANTENNA__1962__A (.DIODE(net610));
 sky130_fd_sc_hd__diode_2 ANTENNA__1963__A (.DIODE(net610));
 sky130_fd_sc_hd__diode_2 ANTENNA__1964__A (.DIODE(net611));
 sky130_fd_sc_hd__diode_2 ANTENNA__1965__A (.DIODE(net611));
 sky130_fd_sc_hd__diode_2 ANTENNA__1966__A (.DIODE(net617));
 sky130_fd_sc_hd__diode_2 ANTENNA__1967__A (.DIODE(net616));
 sky130_fd_sc_hd__diode_2 ANTENNA__1970__A (.DIODE(net616));
 sky130_fd_sc_hd__diode_2 ANTENNA__1971__A (.DIODE(net616));
 sky130_fd_sc_hd__diode_2 ANTENNA__1972__A (.DIODE(net616));
 sky130_fd_sc_hd__diode_2 ANTENNA__1973__A (.DIODE(net616));
 sky130_fd_sc_hd__diode_2 ANTENNA__1974__A (.DIODE(net616));
 sky130_fd_sc_hd__diode_2 ANTENNA__1975__A (.DIODE(net616));
 sky130_fd_sc_hd__diode_2 ANTENNA__1976__A (.DIODE(net616));
 sky130_fd_sc_hd__diode_2 ANTENNA__1977__A (.DIODE(net616));
 sky130_fd_sc_hd__diode_2 ANTENNA__1978__A (.DIODE(net617));
 sky130_fd_sc_hd__diode_2 ANTENNA__1979__A (.DIODE(net616));
 sky130_fd_sc_hd__diode_2 ANTENNA__1995__A (.DIODE(net610));
 sky130_fd_sc_hd__diode_2 ANTENNA__2002__A (.DIODE(net610));
 sky130_fd_sc_hd__diode_2 ANTENNA__2005__A (.DIODE(net609));
 sky130_fd_sc_hd__diode_2 ANTENNA__2007__A (.DIODE(net611));
 sky130_fd_sc_hd__diode_2 ANTENNA__2009__A (.DIODE(net609));
 sky130_fd_sc_hd__diode_2 ANTENNA__2011__A (.DIODE(net609));
 sky130_fd_sc_hd__diode_2 ANTENNA__2016__A (.DIODE(net609));
 sky130_fd_sc_hd__diode_2 ANTENNA__2017__A (.DIODE(net611));
 sky130_fd_sc_hd__diode_2 ANTENNA__2021__A (.DIODE(net609));
 sky130_fd_sc_hd__diode_2 ANTENNA__2022__A (.DIODE(net611));
 sky130_fd_sc_hd__diode_2 ANTENNA__2025__A (.DIODE(net611));
 sky130_fd_sc_hd__diode_2 ANTENNA__2026__A (.DIODE(net611));
 sky130_fd_sc_hd__diode_2 ANTENNA__2027__A (.DIODE(net609));
 sky130_fd_sc_hd__diode_2 ANTENNA__2034__A (.DIODE(net609));
 sky130_fd_sc_hd__diode_2 ANTENNA__2035__A (.DIODE(net612));
 sky130_fd_sc_hd__diode_2 ANTENNA__2036__A (.DIODE(net612));
 sky130_fd_sc_hd__diode_2 ANTENNA__2037__A (.DIODE(net612));
 sky130_fd_sc_hd__diode_2 ANTENNA__2039__A (.DIODE(net617));
 sky130_fd_sc_hd__diode_2 ANTENNA__2040__A (.DIODE(net612));
 sky130_fd_sc_hd__diode_2 ANTENNA__2042__A (.DIODE(net612));
 sky130_fd_sc_hd__diode_2 ANTENNA__2043__A (.DIODE(net612));
 sky130_fd_sc_hd__diode_2 ANTENNA__2044__A (.DIODE(net612));
 sky130_fd_sc_hd__diode_2 ANTENNA__2045__A (.DIODE(net612));
 sky130_fd_sc_hd__diode_2 ANTENNA__2046__A (.DIODE(net612));
 sky130_fd_sc_hd__diode_2 ANTENNA__2047__A (.DIODE(net612));
 sky130_fd_sc_hd__diode_2 ANTENNA__2050__A (.DIODE(net612));
 sky130_fd_sc_hd__diode_2 ANTENNA__2051__A (.DIODE(net612));
 sky130_fd_sc_hd__diode_2 ANTENNA__2053__A (.DIODE(net612));
 sky130_fd_sc_hd__diode_2 ANTENNA__2055__A (.DIODE(net613));
 sky130_fd_sc_hd__diode_2 ANTENNA__2056__A (.DIODE(net613));
 sky130_fd_sc_hd__diode_2 ANTENNA__2057__A (.DIODE(net613));
 sky130_fd_sc_hd__diode_2 ANTENNA__2058__A (.DIODE(net613));
 sky130_fd_sc_hd__diode_2 ANTENNA__2059__A (.DIODE(net613));
 sky130_fd_sc_hd__diode_2 ANTENNA__2060__A (.DIODE(net613));
 sky130_fd_sc_hd__diode_2 ANTENNA__2062__A (.DIODE(net613));
 sky130_fd_sc_hd__diode_2 ANTENNA__2063__A (.DIODE(net613));
 sky130_fd_sc_hd__diode_2 ANTENNA__2064__A (.DIODE(net613));
 sky130_fd_sc_hd__diode_2 ANTENNA__2065__A (.DIODE(net612));
 sky130_fd_sc_hd__diode_2 ANTENNA__2066__A (.DIODE(net613));
 sky130_fd_sc_hd__diode_2 ANTENNA__2067__A (.DIODE(net613));
 sky130_fd_sc_hd__diode_2 ANTENNA__2068__A (.DIODE(net613));
 sky130_fd_sc_hd__diode_2 ANTENNA__2069__A (.DIODE(net613));
 sky130_fd_sc_hd__diode_2 ANTENNA__2161__GATE_N (.DIODE(_0006_));
 sky130_fd_sc_hd__diode_2 ANTENNA_clkbuf_1_0__f_wb_clk_i_A (.DIODE(clknet_0_wb_clk_i));
 sky130_fd_sc_hd__diode_2 ANTENNA_clkbuf_1_1__f_wb_clk_i_A (.DIODE(clknet_0_wb_clk_i));
 sky130_fd_sc_hd__diode_2 ANTENNA_clkbuf_leaf_0_wb_clk_i_A (.DIODE(clknet_1_0__leaf_wb_clk_i));
 sky130_fd_sc_hd__diode_2 ANTENNA_clkbuf_leaf_10_wb_clk_i_A (.DIODE(clknet_1_1__leaf_wb_clk_i));
 sky130_fd_sc_hd__diode_2 ANTENNA_clkbuf_leaf_11_wb_clk_i_A (.DIODE(clknet_1_1__leaf_wb_clk_i));
 sky130_fd_sc_hd__diode_2 ANTENNA_clkbuf_leaf_12_wb_clk_i_A (.DIODE(clknet_1_1__leaf_wb_clk_i));
 sky130_fd_sc_hd__diode_2 ANTENNA_clkbuf_leaf_13_wb_clk_i_A (.DIODE(clknet_1_1__leaf_wb_clk_i));
 sky130_fd_sc_hd__diode_2 ANTENNA_clkbuf_leaf_14_wb_clk_i_A (.DIODE(clknet_1_1__leaf_wb_clk_i));
 sky130_fd_sc_hd__diode_2 ANTENNA_clkbuf_leaf_15_wb_clk_i_A (.DIODE(clknet_1_1__leaf_wb_clk_i));
 sky130_fd_sc_hd__diode_2 ANTENNA_clkbuf_leaf_16_wb_clk_i_A (.DIODE(clknet_1_1__leaf_wb_clk_i));
 sky130_fd_sc_hd__diode_2 ANTENNA_clkbuf_leaf_17_wb_clk_i_A (.DIODE(clknet_1_1__leaf_wb_clk_i));
 sky130_fd_sc_hd__diode_2 ANTENNA_clkbuf_leaf_18_wb_clk_i_A (.DIODE(clknet_1_1__leaf_wb_clk_i));
 sky130_fd_sc_hd__diode_2 ANTENNA_clkbuf_leaf_19_wb_clk_i_A (.DIODE(clknet_1_1__leaf_wb_clk_i));
 sky130_fd_sc_hd__diode_2 ANTENNA_clkbuf_leaf_1_wb_clk_i_A (.DIODE(clknet_1_0__leaf_wb_clk_i));
 sky130_fd_sc_hd__diode_2 ANTENNA_clkbuf_leaf_20_wb_clk_i_A (.DIODE(clknet_1_1__leaf_wb_clk_i));
 sky130_fd_sc_hd__diode_2 ANTENNA_clkbuf_leaf_21_wb_clk_i_A (.DIODE(clknet_1_1__leaf_wb_clk_i));
 sky130_fd_sc_hd__diode_2 ANTENNA_clkbuf_leaf_22_wb_clk_i_A (.DIODE(clknet_1_1__leaf_wb_clk_i));
 sky130_fd_sc_hd__diode_2 ANTENNA_clkbuf_leaf_23_wb_clk_i_A (.DIODE(clknet_1_1__leaf_wb_clk_i));
 sky130_fd_sc_hd__diode_2 ANTENNA_clkbuf_leaf_24_wb_clk_i_A (.DIODE(clknet_1_0__leaf_wb_clk_i));
 sky130_fd_sc_hd__diode_2 ANTENNA_clkbuf_leaf_25_wb_clk_i_A (.DIODE(clknet_1_0__leaf_wb_clk_i));
 sky130_fd_sc_hd__diode_2 ANTENNA_clkbuf_leaf_26_wb_clk_i_A (.DIODE(clknet_1_0__leaf_wb_clk_i));
 sky130_fd_sc_hd__diode_2 ANTENNA_clkbuf_leaf_2_wb_clk_i_A (.DIODE(clknet_1_0__leaf_wb_clk_i));
 sky130_fd_sc_hd__diode_2 ANTENNA_clkbuf_leaf_3_wb_clk_i_A (.DIODE(clknet_1_0__leaf_wb_clk_i));
 sky130_fd_sc_hd__diode_2 ANTENNA_clkbuf_leaf_4_wb_clk_i_A (.DIODE(clknet_1_0__leaf_wb_clk_i));
 sky130_fd_sc_hd__diode_2 ANTENNA_clkbuf_leaf_5_wb_clk_i_A (.DIODE(clknet_1_0__leaf_wb_clk_i));
 sky130_fd_sc_hd__diode_2 ANTENNA_clkbuf_leaf_6_wb_clk_i_A (.DIODE(clknet_1_0__leaf_wb_clk_i));
 sky130_fd_sc_hd__diode_2 ANTENNA_clkbuf_leaf_7_wb_clk_i_A (.DIODE(clknet_1_0__leaf_wb_clk_i));
 sky130_fd_sc_hd__diode_2 ANTENNA_clkbuf_leaf_8_wb_clk_i_A (.DIODE(clknet_1_0__leaf_wb_clk_i));
 sky130_fd_sc_hd__diode_2 ANTENNA_clkbuf_leaf_9_wb_clk_i_A (.DIODE(clknet_1_0__leaf_wb_clk_i));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout521_A (.DIODE(net683));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout522_A (.DIODE(net683));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout523_A (.DIODE(net683));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout524_A (.DIODE(net683));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout525_A (.DIODE(net683));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout527_A (.DIODE(net530));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout528_A (.DIODE(net530));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout529_A (.DIODE(net530));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout531_A (.DIODE(net533));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout532_A (.DIODE(net533));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout534_A (.DIODE(net737));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout536_A (.DIODE(net737));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout537_A (.DIODE(net736));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout538_A (.DIODE(net539));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout539_A (.DIODE(net736));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout540_A (.DIODE(net544));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout542_A (.DIODE(net544));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout543_A (.DIODE(net544));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout544_A (.DIODE(_0946_));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout546_A (.DIODE(net551));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout547_A (.DIODE(net548));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout548_A (.DIODE(net551));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout550_A (.DIODE(net551));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout551_A (.DIODE(_0946_));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout552_A (.DIODE(net555));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout553_A (.DIODE(net555));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout554_A (.DIODE(net555));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout555_A (.DIODE(_0589_));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout556_A (.DIODE(net558));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout557_A (.DIODE(net558));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout558_A (.DIODE(_0589_));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout559_A (.DIODE(_0569_));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout560_A (.DIODE(_0569_));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout561_A (.DIODE(net563));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout562_A (.DIODE(net563));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout563_A (.DIODE(_0569_));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout564_A (.DIODE(net567));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout565_A (.DIODE(net566));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout566_A (.DIODE(net567));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout567_A (.DIODE(_0569_));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout570_A (.DIODE(net571));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout571_A (.DIODE(_0569_));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout572_A (.DIODE(_0007_));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout573_A (.DIODE(_0007_));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout574_A (.DIODE(net576));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout575_A (.DIODE(net576));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout576_A (.DIODE(_0007_));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout577_A (.DIODE(net580));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout578_A (.DIODE(net579));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout579_A (.DIODE(net580));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout580_A (.DIODE(_0007_));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout583_A (.DIODE(net584));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout584_A (.DIODE(_0007_));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout585_A (.DIODE(net588));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout586_A (.DIODE(net588));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout587_A (.DIODE(net588));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout588_A (.DIODE(_0592_));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout589_A (.DIODE(net590));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout590_A (.DIODE(_0592_));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout594_A (.DIODE(_0004_));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout595_A (.DIODE(net597));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout596_A (.DIODE(net597));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout597_A (.DIODE(_0004_));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout598_A (.DIODE(net599));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout599_A (.DIODE(net262));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout600_A (.DIODE(net602));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout601_A (.DIODE(net602));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout602_A (.DIODE(net262));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout603_A (.DIODE(net605));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout604_A (.DIODE(net605));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout605_A (.DIODE(net606));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout606_A (.DIODE(net262));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout607_A (.DIODE(net609));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout608_A (.DIODE(net609));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout609_A (.DIODE(net611));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout610_A (.DIODE(net611));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout611_A (.DIODE(net262));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout615_A (.DIODE(net262));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout616_A (.DIODE(net617));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout617_A (.DIODE(net262));
 sky130_fd_sc_hd__diode_2 ANTENNA_hold113_A (.DIODE(net736));
 sky130_fd_sc_hd__diode_2 ANTENNA_hold127_A (.DIODE(_0796_));
 sky130_fd_sc_hd__diode_2 ANTENNA_hold244_A (.DIODE(_0782_));
 sky130_fd_sc_hd__diode_2 ANTENNA_hold276_A (.DIODE(_0784_));
 sky130_fd_sc_hd__diode_2 ANTENNA_hold298_A (.DIODE(_0690_));
 sky130_fd_sc_hd__diode_2 ANTENNA_hold415_A (.DIODE(_0692_));
 sky130_fd_sc_hd__diode_2 ANTENNA_hold422_A (.DIODE(_0698_));
 sky130_fd_sc_hd__diode_2 ANTENNA_hold443_A (.DIODE(_0696_));
 sky130_fd_sc_hd__diode_2 ANTENNA_hold469_A (.DIODE(net217));
 sky130_fd_sc_hd__diode_2 ANTENNA_hold515_A (.DIODE(_0694_));
 sky130_fd_sc_hd__diode_2 ANTENNA_hold775_A (.DIODE(\reg_temp[98] ));
 sky130_fd_sc_hd__diode_2 ANTENNA_hold786_A (.DIODE(\reg_temp[39] ));
 sky130_fd_sc_hd__diode_2 ANTENNA_hold787_A (.DIODE(\reg_temp[131] ));
 sky130_fd_sc_hd__diode_2 ANTENNA_hold792_A (.DIODE(\reg_temp[46] ));
 sky130_fd_sc_hd__diode_2 ANTENNA_hold793_A (.DIODE(\reg_temp[38] ));
 sky130_fd_sc_hd__diode_2 ANTENNA_hold797_A (.DIODE(\reg_temp[43] ));
 sky130_fd_sc_hd__diode_2 ANTENNA_hold921_A (.DIODE(\reg_temp[32] ));
 sky130_fd_sc_hd__diode_2 ANTENNA_hold922_A (.DIODE(\reg_temp[99] ));
 sky130_fd_sc_hd__diode_2 ANTENNA_hold923_A (.DIODE(\reg_temp[97] ));
 sky130_fd_sc_hd__diode_2 ANTENNA_hold924_A (.DIODE(\reg_temp[143] ));
 sky130_fd_sc_hd__diode_2 ANTENNA_hold925_A (.DIODE(\reg_temp[104] ));
 sky130_fd_sc_hd__diode_2 ANTENNA_hold926_A (.DIODE(\reg_temp[109] ));
 sky130_fd_sc_hd__diode_2 ANTENNA_hold927_A (.DIODE(\reg_temp[24] ));
 sky130_fd_sc_hd__diode_2 ANTENNA_hold929_A (.DIODE(\reg_temp[30] ));
 sky130_fd_sc_hd__diode_2 ANTENNA_hold930_A (.DIODE(\reg_temp[49] ));
 sky130_fd_sc_hd__diode_2 ANTENNA_hold931_A (.DIODE(\reg_temp[126] ));
 sky130_fd_sc_hd__diode_2 ANTENNA_hold932_A (.DIODE(\reg_temp[12] ));
 sky130_fd_sc_hd__diode_2 ANTENNA_hold933_A (.DIODE(\reg_temp[33] ));
 sky130_fd_sc_hd__diode_2 ANTENNA_hold935_A (.DIODE(\reg_temp[116] ));
 sky130_fd_sc_hd__diode_2 ANTENNA_hold937_A (.DIODE(\reg_temp[31] ));
 sky130_fd_sc_hd__diode_2 ANTENNA_hold938_A (.DIODE(\reg_temp[26] ));
 sky130_fd_sc_hd__diode_2 ANTENNA_hold940_A (.DIODE(\reg_temp[34] ));
 sky130_fd_sc_hd__diode_2 ANTENNA_hold941_A (.DIODE(\reg_temp[113] ));
 sky130_fd_sc_hd__diode_2 ANTENNA_hold942_A (.DIODE(\reg_temp[15] ));
 sky130_fd_sc_hd__diode_2 ANTENNA_hold944_A (.DIODE(\reg_temp[112] ));
 sky130_fd_sc_hd__diode_2 ANTENNA_hold945_A (.DIODE(\reg_temp[57] ));
 sky130_fd_sc_hd__diode_2 ANTENNA_hold947_A (.DIODE(\reg_temp[110] ));
 sky130_fd_sc_hd__diode_2 ANTENNA_hold948_A (.DIODE(\reg_temp[120] ));
 sky130_fd_sc_hd__diode_2 ANTENNA_hold949_A (.DIODE(\reg_temp[96] ));
 sky130_fd_sc_hd__diode_2 ANTENNA_hold950_A (.DIODE(\reg_temp[36] ));
 sky130_fd_sc_hd__diode_2 ANTENNA_hold951_A (.DIODE(\reg_temp[4] ));
 sky130_fd_sc_hd__diode_2 ANTENNA_hold953_A (.DIODE(\reg_temp[95] ));
 sky130_fd_sc_hd__diode_2 ANTENNA_hold955_A (.DIODE(\reg_temp[103] ));
 sky130_fd_sc_hd__diode_2 ANTENNA_hold956_A (.DIODE(\reg_temp[27] ));
 sky130_fd_sc_hd__diode_2 ANTENNA_hold957_A (.DIODE(\reg_temp[138] ));
 sky130_fd_sc_hd__diode_2 ANTENNA_hold958_A (.DIODE(\reg_temp[5] ));
 sky130_fd_sc_hd__diode_2 ANTENNA_hold959_A (.DIODE(\reg_temp[114] ));
 sky130_fd_sc_hd__diode_2 ANTENNA_hold95_A (.DIODE(_0750_));
 sky130_fd_sc_hd__diode_2 ANTENNA_hold961_A (.DIODE(\reg_temp[121] ));
 sky130_fd_sc_hd__diode_2 ANTENNA_hold962_A (.DIODE(\reg_temp[28] ));
 sky130_fd_sc_hd__diode_2 ANTENNA_hold963_A (.DIODE(\reg_temp[18] ));
 sky130_fd_sc_hd__diode_2 ANTENNA_hold964_A (.DIODE(\reg_temp[19] ));
 sky130_fd_sc_hd__diode_2 ANTENNA_hold965_A (.DIODE(\reg_temp[3] ));
 sky130_fd_sc_hd__diode_2 ANTENNA_hold966_A (.DIODE(\reg_temp[101] ));
 sky130_fd_sc_hd__diode_2 ANTENNA_hold967_A (.DIODE(\reg_temp[87] ));
 sky130_fd_sc_hd__diode_2 ANTENNA_hold968_A (.DIODE(\reg_temp[119] ));
 sky130_fd_sc_hd__diode_2 ANTENNA_hold969_A (.DIODE(\reg_temp[25] ));
 sky130_fd_sc_hd__diode_2 ANTENNA_hold970_A (.DIODE(\reg_temp[100] ));
 sky130_fd_sc_hd__diode_2 ANTENNA_hold971_A (.DIODE(\reg_temp[82] ));
 sky130_fd_sc_hd__diode_2 ANTENNA_hold972_A (.DIODE(\reg_temp[13] ));
 sky130_fd_sc_hd__diode_2 ANTENNA_hold973_A (.DIODE(\reg_temp[21] ));
 sky130_fd_sc_hd__diode_2 ANTENNA_hold974_A (.DIODE(\reg_temp[139] ));
 sky130_fd_sc_hd__diode_2 ANTENNA_hold975_A (.DIODE(\reg_temp[102] ));
 sky130_fd_sc_hd__diode_2 ANTENNA_hold976_A (.DIODE(\reg_temp[123] ));
 sky130_fd_sc_hd__diode_2 ANTENNA_hold977_A (.DIODE(\reg_temp[89] ));
 sky130_fd_sc_hd__diode_2 ANTENNA_hold978_A (.DIODE(\reg_temp[115] ));
 sky130_fd_sc_hd__diode_2 ANTENNA_hold979_A (.DIODE(\reg_temp[86] ));
 sky130_fd_sc_hd__diode_2 ANTENNA_hold980_A (.DIODE(\reg_temp[20] ));
 sky130_fd_sc_hd__diode_2 ANTENNA_hold981_A (.DIODE(\reg_temp[22] ));
 sky130_fd_sc_hd__diode_2 ANTENNA_hold982_A (.DIODE(\reg_temp[29] ));
 sky130_fd_sc_hd__diode_2 ANTENNA_hold983_A (.DIODE(\reg_temp[4] ));
 sky130_fd_sc_hd__diode_2 ANTENNA_hold984_A (.DIODE(\reg_temp[85] ));
 sky130_fd_sc_hd__diode_2 ANTENNA_hold985_A (.DIODE(\reg_temp[17] ));
 sky130_fd_sc_hd__diode_2 ANTENNA_hold986_A (.DIODE(\reg_temp[105] ));
 sky130_fd_sc_hd__diode_2 ANTENNA_hold987_A (.DIODE(\reg_temp[35] ));
 sky130_fd_sc_hd__diode_2 ANTENNA_hold988_A (.DIODE(\reg_temp[92] ));
 sky130_fd_sc_hd__diode_2 ANTENNA_hold989_A (.DIODE(\reg_temp[41] ));
 sky130_fd_sc_hd__diode_2 ANTENNA_hold990_A (.DIODE(\reg_temp[23] ));
 sky130_fd_sc_hd__diode_2 ANTENNA_hold991_A (.DIODE(\reg_temp[40] ));
 sky130_fd_sc_hd__diode_2 ANTENNA_hold992_A (.DIODE(\reg_temp[93] ));
 sky130_fd_sc_hd__diode_2 ANTENNA_hold993_A (.DIODE(\reg_temp[8] ));
 sky130_fd_sc_hd__diode_2 ANTENNA_output263_A (.DIODE(net263));
 sky130_fd_sc_hd__diode_2 ANTENNA_output288_A (.DIODE(net288));
 sky130_fd_sc_hd__diode_2 ANTENNA_output292_A (.DIODE(net292));
 sky130_fd_sc_hd__diode_2 ANTENNA_output361_A (.DIODE(net361));
 sky130_fd_sc_hd__diode_2 ANTENNA_output365_A (.DIODE(net365));
 sky130_fd_sc_hd__diode_2 ANTENNA_output402_A (.DIODE(net402));
 sky130_fd_sc_hd__diode_2 ANTENNA_output405_A (.DIODE(net405));
 sky130_fd_sc_hd__diode_2 ANTENNA_output406_A (.DIODE(net406));
 sky130_fd_sc_hd__diode_2 ANTENNA_output407_A (.DIODE(net407));
 sky130_fd_sc_hd__diode_2 ANTENNA_output451_A (.DIODE(net1285));
 sky130_fd_sc_hd__diode_2 ANTENNA_output453_A (.DIODE(net1315));
 sky130_fd_sc_hd__diode_2 ANTENNA_output465_A (.DIODE(net1227));
 sky130_fd_sc_hd__diode_2 ANTENNA_output475_A (.DIODE(net1225));
 sky130_fd_sc_hd__diode_2 ANTENNA_output480_A (.DIODE(net1304));
 sky130_fd_sc_hd__diode_2 ANTENNA_output484_A (.DIODE(net1303));
 sky130_fd_sc_hd__fill_1 FILLER_0_0_141 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_0_253 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_0_298 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_0_3 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_0_365 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_0_369 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_0_391 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_0_402 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_0_424 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_0_559 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_0_573 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_0_592 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_0_612 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_0_615 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_0_62 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_0_642 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_0_699 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_0_712 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_0_80 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_10_128 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_10_138 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_10_219 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_10_222 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_10_233 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_10_250 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_10_264 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_10_290 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_10_3 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_10_305 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_10_309 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_10_315 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_10_342 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_10_345 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_10_348 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_10_372 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_10_415 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_10_418 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_10_433 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_10_475 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_10_513 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_10_531 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_10_584 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_10_587 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_10_651 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_10_699 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_10_701 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_10_713 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_11_135 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_11_143 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_11_20 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_11_214 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_11_228 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_11_238 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_11_258 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_11_270 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_11_298 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_11_3 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_11_310 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_11_333 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_11_348 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_11_383 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_11_400 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_11_410 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_11_419 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_11_422 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_11_447 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_11_497 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_11_501 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_11_505 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_11_509 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_11_558 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_11_583 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_11_628 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_12_11 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_12_158 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_12_171 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_12_197 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_12_213 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_12_230 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_12_233 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_12_250 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_12_253 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_12_290 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_12_3 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_12_301 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_12_307 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_12_309 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_12_341 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_12_344 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_12_35 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_12_356 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_12_371 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_12_374 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_12_38 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_12_387 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_12_419 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_12_424 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_12_432 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_12_436 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_12_439 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_12_442 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_12_447 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_12_508 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_12_527 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_12_530 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_12_55 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_12_58 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_12_581 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_12_61 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_12_661 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_12_690 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_12_71 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_12_713 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_12_8 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_12_80 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_12_93 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_13_174 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_13_183 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_13_22 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_13_225 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_13_238 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_13_245 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_13_257 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_13_269 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_13_276 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_13_281 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_13_288 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_13_300 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_13_326 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_13_331 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_13_334 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_13_337 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_13_345 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_13_353 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_13_361 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_13_366 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_13_372 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_13_376 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_13_388 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_13_393 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_13_405 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_13_426 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_13_438 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_13_449 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_13_452 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_13_496 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_13_499 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_13_503 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_13_515 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_13_63 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_13_637 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_13_661 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_13_688 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_13_691 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_13_700 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_13_711 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_14_14 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_14_163 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_14_175 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_14_183 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_14_187 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_14_197 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_14_20 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_14_205 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_14_214 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_14_222 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_14_226 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_14_229 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_14_241 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_14_249 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_14_253 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_14_265 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_14_277 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_14_289 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_14_29 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_14_3 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_14_301 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_14_307 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_14_309 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_14_313 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_14_316 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_14_328 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_14_340 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_14_352 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_14_376 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_14_379 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_14_391 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_14_403 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_14_421 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_14_445 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_14_451 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_14_454 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_14_469 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_14_475 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_14_477 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_14_485 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_14_516 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_14_533 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_14_542 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_14_587 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_14_610 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_14_619 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_14_622 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_14_642 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_14_653 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_14_662 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_14_666 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_14_669 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_14_672 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_14_675 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_14_678 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_14_699 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_14_701 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_14_85 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_14_99 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_15_113 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_15_136 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_15_15 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_15_158 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_15_192 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_15_199 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_15_20 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_15_215 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_15_218 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_15_221 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_15_225 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_15_23 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_15_237 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_15_249 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_15_259 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_15_271 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_15_279 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_15_281 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_15_293 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_15_3 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_15_301 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_15_319 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_15_323 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_15_326 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_15_334 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_15_337 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_15_343 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_15_369 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_15_376 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_15_379 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_15_391 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_15_393 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_15_405 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_15_411 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_15_414 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_15_426 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_15_438 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_15_446 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_15_449 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_15_461 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_15_473 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_15_481 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_15_49 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_15_491 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_15_505 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_15_524 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_15_527 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_15_564 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_15_57 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_15_608 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_15_612 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_15_615 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_15_617 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_15_620 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_15_623 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_15_626 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_15_635 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_15_638 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_15_64 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_15_641 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_15_644 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_15_647 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_15_656 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_15_659 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_15_662 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_15_665 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_15_668 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_15_67 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_15_671 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_15_681 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_15_689 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_15_708 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_15_92 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_16_10 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_16_102 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_16_127 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_16_13 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_16_136 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_16_16 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_16_19 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_16_193 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_16_197 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_16_200 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_16_203 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_16_214 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_16_217 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_16_229 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_16_241 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_16_249 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_16_256 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_16_268 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_16_271 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_16_283 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_16_286 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_16_298 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_16_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_16_332 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_16_344 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_16_362 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_16_365 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_16_376 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_16_388 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_16_400 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_16_404 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_16_408 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_16_413 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_16_416 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_16_419 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_16_428 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_16_432 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_16_444 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_16_456 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_16_468 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_16_477 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_16_489 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_16_510 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_16_52 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_16_521 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_16_533 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_16_565 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_16_568 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_16_57 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_16_571 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_16_582 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_16_586 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_16_589 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_16_626 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_16_629 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_16_63 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_16_632 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_16_635 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_16_638 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_16_641 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_16_645 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_16_648 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_16_651 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_16_654 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_16_657 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_16_660 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_16_672 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_16_684 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_16_694 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_16_697 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_16_7 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_16_701 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_16_704 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_16_707 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_16_713 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_16_82 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_16_85 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_17_104 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_17_110 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_17_12 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_17_124 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_17_128 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_17_142 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_17_15 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_17_164 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_17_197 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_17_200 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_17_212 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_17_222 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_17_225 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_17_237 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_17_251 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_17_255 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_17_259 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_17_262 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_17_265 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_17_274 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_17_279 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_17_284 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_17_287 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_17_296 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_17_3 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_17_310 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_17_326 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_17_334 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_17_337 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_17_343 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_17_355 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_17_358 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_17_363 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_17_378 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_17_393 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_17_41 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_17_415 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_17_438 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_17_442 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_17_45 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_17_457 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_17_478 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_17_483 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_17_488 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_17_498 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_17_501 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_17_505 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_17_517 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_17_523 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_17_526 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_17_529 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_17_55 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_17_552 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_17_564 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_17_567 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_17_57 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_17_570 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_17_573 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_17_576 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_17_579 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_17_595 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_17_6 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_17_60 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_17_617 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_17_63 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_17_637 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_17_661 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_17_669 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_17_673 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_17_685 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_17_697 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_17_709 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_17_713 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_17_85 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_17_9 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_18_10 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_18_103 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_18_123 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_18_13 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_18_138 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_18_16 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_18_164 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_18_193 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_18_205 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_18_211 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_18_230 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_18_233 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_18_236 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_18_242 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_18_245 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_18_251 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_18_262 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_18_29 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_18_297 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_18_3 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_18_305 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_18_309 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_18_314 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_18_318 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_18_327 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_18_339 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_18_343 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_18_346 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_18_361 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_18_365 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_18_368 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_18_372 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_18_378 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_18_389 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_18_399 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_18_447 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_18_47 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_18_474 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_18_477 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_18_480 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_18_50 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_18_501 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_18_504 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_18_508 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_18_511 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_18_523 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_18_53 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_18_531 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_18_540 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_18_546 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_18_568 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_18_571 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_18_575 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_18_578 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_18_583 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_18_589 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_18_596 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_18_600 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_18_603 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_18_633 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_18_643 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_18_653 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_18_656 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_18_659 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_18_663 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_18_687 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_18_699 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_18_7 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_18_701 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_18_713 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_18_96 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_19_103 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_19_11 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_19_127 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_19_152 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_19_155 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_19_160 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_19_164 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_19_167 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_19_169 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_19_172 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_19_201 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_19_208 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_19_220 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_19_225 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_19_234 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_19_237 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_19_278 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_19_3 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_19_301 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_19_309 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_19_317 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_19_326 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_19_329 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_19_335 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_19_337 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_19_346 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_19_363 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_19_378 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_19_381 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_19_384 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_19_390 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_19_413 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_19_422 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_19_426 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_19_447 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_19_449 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_19_463 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_19_466 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_19_486 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_19_489 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_19_500 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_19_503 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_19_519 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_19_522 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_19_53 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_19_535 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_19_538 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_19_542 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_19_545 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_19_551 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_19_554 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_19_561 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_19_57 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_19_573 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_19_581 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_19_585 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_19_589 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_19_593 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_19_596 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_19_599 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_19_604 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_19_62 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_19_625 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_19_637 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_19_648 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_19_65 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_19_651 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_19_655 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_19_666 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_19_673 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_19_685 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_19_697 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_19_7 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_19_709 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_19_713 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_1_220 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_1_223 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_1_281 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_1_330 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_1_342 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_1_354 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_1_366 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_1_378 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_1_385 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_1_389 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_1_411 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_1_444 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_1_670 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_1_68 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_1_681 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_1_79 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_20_120 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_20_127 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_20_141 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_20_15 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_20_153 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_20_157 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_20_160 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_20_173 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_20_177 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_20_188 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_20_195 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_20_197 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_20_204 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_20_207 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_20_219 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_20_23 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_20_231 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_20_243 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_20_249 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_20_256 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_20_261 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_20_264 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_20_298 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_20_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_20_317 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_20_329 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_20_341 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_20_345 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_20_348 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_20_356 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_20_359 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_20_362 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_20_365 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_20_37 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_20_394 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_20_40 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_20_402 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_20_405 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_20_408 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_20_414 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_20_421 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_20_433 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_20_44 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_20_47 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_20_473 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_20_477 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_20_489 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_20_494 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_20_503 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_20_506 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_20_512 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_20_528 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_20_53 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_20_531 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_20_533 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_20_536 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_20_539 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_20_547 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_20_551 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_20_56 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_20_580 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_20_589 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_20_59 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_20_601 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_20_607 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_20_629 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_20_632 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_20_687 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_20_699 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_20_701 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_20_713 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_20_80 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_20_85 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_21_103 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_21_106 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_21_109 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_21_124 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_21_127 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_21_130 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_21_134 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_21_137 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_21_147 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_21_15 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_21_151 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_21_154 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_21_157 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_21_160 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_21_169 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_21_181 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_21_187 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_21_199 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_21_216 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_21_219 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_21_223 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_21_225 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_21_229 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_21_23 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_21_235 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_21_247 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_21_255 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_21_260 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_21_266 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_21_276 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_21_279 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_21_281 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_21_294 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_21_297 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_21_3 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_21_309 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_21_317 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_21_323 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_21_335 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_21_337 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_21_345 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_21_352 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_21_36 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_21_373 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_21_386 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_21_389 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_21_409 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_21_426 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_21_434 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_21_437 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_21_444 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_21_447 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_21_449 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_21_455 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_21_461 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_21_464 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_21_467 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_21_470 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_21_48 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_21_482 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_21_486 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_21_489 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_21_500 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_21_505 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_21_517 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_21_57 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_21_581 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_21_609 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_21_612 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_21_617 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_21_621 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_21_630 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_21_642 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_21_662 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_21_665 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_21_671 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_21_673 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_21_681 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_21_702 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_21_80 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_21_83 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_21_86 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_21_98 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_22_129 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_22_133 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_22_137 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_22_149 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_22_15 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_22_161 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_22_165 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_22_168 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_22_179 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_22_191 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_22_207 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_22_214 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_22_238 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_22_250 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_22_253 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_22_261 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_22_265 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_22_268 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_22_27 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_22_29 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_22_296 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_22_299 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_22_3 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_22_307 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_22_309 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_22_321 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_22_333 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_22_340 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_22_344 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_22_347 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_22_365 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_22_390 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_22_402 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_22_414 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_22_421 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_22_433 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_22_439 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_22_447 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_22_450 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_22_462 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_22_466 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_22_474 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_22_477 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_22_485 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_22_488 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_22_49 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_22_518 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_22_52 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_22_527 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_22_539 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_22_549 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_22_553 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_22_597 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_22_604 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_22_607 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_22_613 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_22_625 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_22_637 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_22_64 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_22_641 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_22_665 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_22_673 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_22_709 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_22_713 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_22_76 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_22_85 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_22_91 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_22_94 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_23_103 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_23_11 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_23_110 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_23_113 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_23_123 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_23_126 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_23_129 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_23_132 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_23_135 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_23_147 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_23_161 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_23_165 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_23_169 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_23_189 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_23_192 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_23_195 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_23_223 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_23_236 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_23_239 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_23_260 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_23_266 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_23_269 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_23_277 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_23_292 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_23_295 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_23_298 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_23_3 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_23_301 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_23_309 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_23_321 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_23_324 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_23_337 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_23_353 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_23_357 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_23_362 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_23_365 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_23_37 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_23_375 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_23_384 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_23_409 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_23_421 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_23_427 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_23_439 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_23_443 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_23_449 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_23_454 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_23_457 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_23_460 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_23_474 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_23_477 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_23_481 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_23_484 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_23_487 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_23_49 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_23_499 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_23_503 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_23_505 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_23_511 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_23_521 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_23_530 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_23_536 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_23_541 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_23_544 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_23_547 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_23_556 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_23_561 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_23_596 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_23_606 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_23_614 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_23_617 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_23_629 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_23_637 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_23_644 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_23_670 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_23_700 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_23_712 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_23_80 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_23_92 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_24_101 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_24_107 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_24_121 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_24_141 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_24_15 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_24_159 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_24_163 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_24_167 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_24_19 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_24_192 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_24_197 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_24_209 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_24_233 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_24_241 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_24_246 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_24_249 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_24_253 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_24_26 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_24_3 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_24_301 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_24_304 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_24_332 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_24_344 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_24_356 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_24_37 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_24_374 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_24_377 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_24_380 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_24_391 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_24_394 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_24_402 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_24_405 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_24_408 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_24_417 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_24_441 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_24_45 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_24_462 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_24_471 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_24_48 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_24_480 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_24_483 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_24_494 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_24_502 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_24_505 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_24_509 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_24_523 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_24_531 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_24_533 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_24_545 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_24_575 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_24_587 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_24_589 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_24_601 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_24_613 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_24_625 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_24_637 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_24_643 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_24_645 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_24_657 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_24_662 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_24_668 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_24_677 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_24_687 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_24_690 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_24_693 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_24_699 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_24_701 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_24_713 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_24_73 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_24_76 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_24_79 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_24_83 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_24_85 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_24_97 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_25_110 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_25_113 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_25_116 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_25_128 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_25_163 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_25_167 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_25_192 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_25_213 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_25_234 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_25_237 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_25_240 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_25_246 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_25_270 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_25_3 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_25_333 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_25_337 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_25_349 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_25_361 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_25_373 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_25_377 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_25_380 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_25_383 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_25_386 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_25_393 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_25_401 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_25_408 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_25_412 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_25_417 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_25_43 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_25_486 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_25_496 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_25_499 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_25_502 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_25_525 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_25_528 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_25_532 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_25_538 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_25_542 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_25_545 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_25_557 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_25_561 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_25_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_25_573 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_25_585 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_25_593 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_25_597 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_25_603 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_25_615 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_25_617 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_25_625 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_25_628 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_25_631 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_25_643 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_25_655 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_25_667 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_25_671 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_25_673 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_25_682 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_25_694 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_25_706 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_25_78 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_25_81 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_25_84 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_25_96 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_26_128 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_26_136 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_26_141 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_26_15 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_26_156 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_26_165 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_26_170 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_26_191 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_26_197 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_26_208 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_26_222 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_26_225 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_26_232 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_26_244 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_26_253 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_26_264 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_26_269 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_26_27 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_26_272 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_26_275 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_26_29 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_26_294 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_26_297 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_26_3 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_26_326 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_26_329 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_26_33 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_26_341 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_26_353 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_26_361 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_26_365 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_26_370 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_26_373 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_26_376 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_26_386 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_26_392 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_26_395 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_26_41 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_26_416 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_26_421 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_26_425 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_26_438 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_26_448 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_26_451 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_26_472 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_26_475 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_26_477 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_26_481 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_26_512 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_26_515 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_26_518 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_26_530 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_26_553 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_26_556 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_26_568 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_26_580 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_26_589 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_26_613 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_26_616 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_26_640 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_26_645 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_26_654 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_26_658 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_26_661 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_26_673 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_26_685 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_26_697 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_26_701 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_26_713 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_26_74 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_26_82 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_26_85 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_27_103 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_27_113 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_27_116 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_27_15 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_27_150 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_27_154 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_27_157 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_27_165 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_27_169 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_27_173 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_27_188 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_27_193 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_27_196 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_27_199 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_27_205 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_27_209 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_27_219 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_27_222 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_27_23 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_27_248 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_27_252 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_27_261 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_27_266 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_27_278 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_27_281 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_27_294 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_27_3 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_27_303 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_27_306 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_27_316 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_27_328 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_27_337 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_27_349 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_27_355 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_27_363 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_27_381 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_27_390 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_27_393 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_27_401 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_27_409 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_27_41 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_27_445 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_27_455 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_27_458 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_27_47 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_27_473 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_27_481 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_27_503 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_27_509 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_27_512 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_27_521 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_27_534 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_27_537 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_27_558 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_27_569 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_27_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_27_581 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_27_593 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_27_615 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_27_620 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_27_670 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_27_673 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_27_679 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_27_68 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_27_703 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_27_711 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_27_72 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_27_75 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_27_87 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_27_99 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_28_105 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_28_110 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_28_113 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_28_116 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_28_15 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_28_152 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_28_155 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_28_158 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_28_193 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_28_197 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_28_205 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_28_208 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_28_211 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_28_214 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_28_217 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_28_240 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_28_243 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_28_246 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_28_253 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_28_261 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_28_265 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_28_27 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_28_277 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_28_283 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_28_286 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_28_289 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_28_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_28_295 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_28_3 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_28_307 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_28_309 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_28_312 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_28_344 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_28_347 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_28_351 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_28_355 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_28_363 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_28_365 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_28_39 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_28_398 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_28_410 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_28_418 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_28_421 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_28_426 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_28_429 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_28_450 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_28_455 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_28_458 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_28_461 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_28_464 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_28_473 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_28_477 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_28_489 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_28_497 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_28_51 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_28_516 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_28_525 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_28_528 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_28_531 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_28_533 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_28_536 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_28_557 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_28_561 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_28_57 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_28_582 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_28_586 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_28_589 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_28_636 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_28_662 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_28_674 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_28_696 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_28_701 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_28_71 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_28_713 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_28_74 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_28_82 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_28_85 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_28_97 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_29_111 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_29_121 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_29_124 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_29_132 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_29_146 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_29_15 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_29_162 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_29_169 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_29_172 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_29_183 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_29_206 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_29_219 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_29_222 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_29_237 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_29_240 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_29_243 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_29_253 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_29_27 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_29_277 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_29_281 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_29_289 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_29_294 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_29_297 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_29_3 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_29_308 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_29_330 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_29_333 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_29_337 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_29_349 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_29_373 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_29_379 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_29_382 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_29_385 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_29_389 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_29_393 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_29_396 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_29_406 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_29_41 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_29_427 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_29_435 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_29_44 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_29_443 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_29_446 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_29_466 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_29_469 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_29_477 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_29_482 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_29_485 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_29_489 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_29_501 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_29_505 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_29_508 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_29_511 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_29_514 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_29_541 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_29_544 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_29_547 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_29_554 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_29_57 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_29_577 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_29_607 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_29_61 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_29_610 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_29_613 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_29_617 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_29_629 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_29_643 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_29_65 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_29_654 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_29_668 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_29_673 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_29_679 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_29_69 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_29_691 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_29_703 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_29_711 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_29_78 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_29_90 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_2_104 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_2_141 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_2_165 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_2_197 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_2_216 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_2_219 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_2_253 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_2_264 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_2_289 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_2_306 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_2_328 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_2_334 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_2_341 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_2_347 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_2_359 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_2_363 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_2_365 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_2_377 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_2_389 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_2_401 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_2_405 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_2_418 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_2_448 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_2_565 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_2_57 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_2_586 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_2_592 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_2_699 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_2_701 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_2_713 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_2_93 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_30_122 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_30_125 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_30_129 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_30_141 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_30_145 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_30_148 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_30_15 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_30_155 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_30_167 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_30_178 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_30_190 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_30_193 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_30_197 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_30_200 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_30_21 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_30_242 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_30_246 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_30_25 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_30_253 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_30_286 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_30_29 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_30_298 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_30_3 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_30_309 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_30_354 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_30_382 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_30_385 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_30_393 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_30_397 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_30_409 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_30_421 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_30_43 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_30_438 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_30_454 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_30_457 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_30_469 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_30_473 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_30_495 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_30_499 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_30_502 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_30_505 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_30_508 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_30_512 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_30_515 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_30_531 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_30_547 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_30_550 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_30_553 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_30_557 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_30_560 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_30_563 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_30_572 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_30_580 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_30_587 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_30_589 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_30_599 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_30_609 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_30_621 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_30_633 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_30_641 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_30_645 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_30_657 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_30_660 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_30_672 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_30_678 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_30_699 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_30_704 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_30_707 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_30_713 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_30_74 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_30_82 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_30_85 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_30_89 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_31_11 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_31_125 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_31_128 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_31_162 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_31_165 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_31_169 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_31_183 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_31_189 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_31_210 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_31_234 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_31_237 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_31_249 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_31_253 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_31_279 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_31_290 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_31_293 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_31_3 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_31_304 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_31_315 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_31_318 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_31_327 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_31_330 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_31_345 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_31_357 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_31_371 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_31_374 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_31_377 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_31_387 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_31_391 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_31_393 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_31_398 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_31_401 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_31_410 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_31_430 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_31_442 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_31_445 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_31_449 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_31_45 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_31_459 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_31_462 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_31_472 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_31_475 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_31_484 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_31_487 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_31_492 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_31_503 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_31_512 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_31_52 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_31_544 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_31_547 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_31_550 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_31_558 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_31_561 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_31_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_31_573 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_31_585 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_31_597 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_31_609 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_31_615 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_31_617 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_31_629 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_31_641 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_31_653 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_31_665 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_31_671 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_31_673 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_31_704 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_31_707 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_31_713 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_31_76 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_31_79 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_31_82 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_31_88 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_32_126 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_32_129 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_32_150 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_32_154 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_32_157 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_32_194 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_32_197 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_32_203 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_32_227 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_32_230 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_32_242 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_32_253 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_32_256 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_32_292 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_32_3 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_32_300 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_32_305 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_32_309 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_32_319 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_32_32 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_32_327 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_32_353 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_32_361 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_32_365 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_32_373 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_32_377 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_32_384 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_32_387 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_32_390 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_32_400 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_32_404 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_32_408 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_32_411 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_32_419 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_32_421 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_32_433 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_32_441 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_32_464 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_32_497 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_32_518 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_32_540 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_32_557 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_32_576 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_32_589 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_32_596 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_32_599 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_32_604 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_32_611 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_32_614 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_32_622 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_32_637 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_32_643 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_32_645 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_32_657 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_32_668 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_32_671 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_32_694 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_32_709 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_32_712 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_32_82 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_32_85 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_33_107 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_33_111 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_33_113 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_33_118 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_33_121 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_33_133 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_33_140 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_33_15 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_33_150 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_33_153 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_33_165 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_33_169 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_33_183 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_33_186 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_33_198 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_33_206 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_33_221 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_33_239 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_33_242 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_33_254 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_33_262 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_33_267 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_33_279 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_33_281 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_33_284 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_33_292 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_33_3 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_33_317 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_33_33 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_33_330 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_33_333 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_33_345 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_33_357 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_33_365 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_33_370 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_33_378 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_33_386 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_33_389 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_33_393 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_33_414 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_33_422 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_33_427 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_33_43 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_33_430 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_33_438 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_33_442 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_33_457 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_33_462 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_33_474 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_33_477 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_33_500 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_33_503 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_33_544 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_33_547 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_33_57 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_33_581 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_33_585 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_33_593 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_33_612 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_33_643 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_33_651 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_33_681 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_33_701 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_33_707 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_33_710 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_33_713 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_33_83 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_33_86 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_33_98 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_34_105 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_34_117 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_34_129 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_34_137 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_34_141 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_34_15 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_34_154 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_34_162 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_34_187 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_34_195 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_34_197 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_34_203 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_34_222 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_34_23 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_34_236 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_34_249 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_34_253 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_34_265 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_34_270 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_34_278 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_34_281 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_34_287 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_34_290 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_34_294 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_34_297 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_34_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_34_320 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_34_332 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_34_344 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_34_356 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_34_360 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_34_363 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_34_37 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_34_370 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_34_373 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_34_387 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_34_390 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_34_399 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_34_402 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_34_405 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_34_413 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_34_416 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_34_45 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_34_454 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_34_462 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_34_465 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_34_475 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_34_477 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_34_480 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_34_501 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_34_510 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_34_520 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_34_531 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_34_533 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_34_541 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_34_547 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_34_567 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_34_571 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_34_580 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_34_583 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_34_587 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_34_589 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_34_597 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_34_610 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_34_62 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_34_636 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_34_66 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_34_662 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_34_665 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_34_673 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_34_685 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_34_699 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_34_701 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_34_705 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_34_708 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_34_71 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_34_711 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_34_74 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_34_83 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_34_85 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_34_93 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_35_103 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_35_111 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_35_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_35_118 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_35_130 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_35_15 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_35_156 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_35_159 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_35_162 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_35_169 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_35_189 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_35_192 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_35_198 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_35_222 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_35_225 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_35_228 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_35_231 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_35_258 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_35_266 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_35_293 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_35_297 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_35_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_35_309 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_35_321 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_35_325 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_35_329 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_35_335 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_35_337 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_35_349 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_35_361 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_35_373 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_35_377 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_35_380 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_35_387 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_35_390 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_35_40 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_35_402 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_35_405 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_35_409 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_35_427 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_35_430 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_35_433 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_35_442 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_35_449 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_35_45 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_35_452 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_35_473 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_35_485 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_35_497 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_35_501 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_35_508 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_35_511 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_35_514 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_35_517 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_35_525 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_35_535 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_35_547 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_35_557 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_35_57 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_35_572 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_35_575 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_35_587 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_35_599 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_35_605 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_35_614 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_35_617 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_35_622 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_35_628 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_35_631 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_35_643 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_35_66 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_35_665 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_35_671 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_35_673 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_35_685 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_35_689 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_35_69 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_35_695 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_35_700 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_35_703 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_35_706 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_35_709 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_35_712 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_36_104 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_36_128 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_36_136 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_36_15 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_36_163 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_36_167 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_36_186 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_36_189 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_36_195 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_36_197 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_36_224 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_36_247 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_36_251 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_36_261 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_36_264 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_36_27 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_36_291 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_36_3 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_36_309 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_36_360 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_36_373 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_36_378 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_36_399 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_36_40 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_36_411 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_36_415 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_36_418 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_36_421 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_36_433 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_36_445 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_36_451 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_36_458 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_36_461 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_36_469 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_36_472 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_36_475 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_36_486 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_36_498 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_36_510 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_36_516 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_36_519 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_36_530 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_36_544 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_36_547 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_36_559 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_36_571 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_36_583 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_36_587 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_36_594 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_36_597 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_36_605 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_36_615 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_36_623 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_36_627 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_36_63 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_36_635 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_36_645 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_36_66 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_36_661 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_36_669 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_36_673 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_36_677 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_36_698 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_36_701 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_36_704 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_36_707 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_36_710 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_36_713 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_36_78 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_36_83 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_37_109 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_37_122 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_37_128 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_37_15 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_37_162 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_37_169 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_37_178 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_37_191 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_37_194 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_37_222 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_37_225 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_37_228 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_37_234 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_37_251 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_37_254 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_37_262 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_37_27 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_37_275 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_37_278 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_37_281 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_37_3 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_37_301 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_37_304 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_37_308 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_37_311 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_37_33 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_37_331 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_37_354 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_37_366 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_37_393 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_37_396 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_37_399 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_37_411 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_37_416 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_37_419 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_37_430 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_37_442 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_37_449 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_37_461 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_37_473 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_37_485 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_37_497 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_37_503 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_37_505 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_37_51 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_37_517 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_37_536 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_37_539 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_37_55 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_37_551 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_37_559 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_37_561 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_37_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_37_573 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_37_585 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_37_597 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_37_60 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_37_609 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_37_615 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_37_617 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_37_623 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_37_626 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_37_655 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_37_661 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_37_670 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_37_673 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_37_676 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_37_68 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_37_680 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_37_691 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_37_694 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_37_697 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_37_700 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_37_709 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_37_712 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_38_102 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_38_105 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_38_108 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_38_127 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_38_137 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_38_15 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_38_157 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_38_160 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_38_189 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_38_192 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_38_197 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_38_209 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_38_213 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_38_217 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_38_220 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_38_228 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_38_256 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_38_259 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_38_267 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_38_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_38_272 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_38_284 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_38_29 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_38_292 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_38_295 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_38_3 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_38_307 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_38_309 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_38_317 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_38_320 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_38_324 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_38_33 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_38_336 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_38_348 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_38_360 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_38_365 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_38_375 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_38_378 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_38_394 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_38_405 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_38_41 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_38_417 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_38_421 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_38_429 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_38_437 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_38_449 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_38_45 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_38_460 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_38_463 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_38_475 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_38_477 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_38_489 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_38_501 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_38_509 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_38_514 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_38_519 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_38_522 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_38_530 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_38_533 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_38_545 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_38_557 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_38_561 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_38_57 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_38_571 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_38_574 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_38_580 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_38_583 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_38_587 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_38_598 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_38_617 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_38_629 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_38_653 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_38_658 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_38_661 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_38_664 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_38_667 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_38_670 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_38_673 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_38_677 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_38_680 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_38_683 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_38_686 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_38_689 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_38_69 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_38_704 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_38_75 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_39_101 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_39_104 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_39_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_39_121 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_39_133 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_39_145 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_39_15 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_39_151 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_39_163 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_39_167 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_39_169 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_39_207 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_39_219 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_39_223 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_39_225 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_39_247 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_39_250 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_39_262 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_39_274 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_39_281 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_39_285 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_39_297 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_39_3 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_39_301 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_39_304 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_39_315 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_39_332 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_39_337 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_39_349 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_39_375 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_39_378 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_39_381 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_39_389 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_39_399 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_39_402 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_39_410 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_39_422 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_39_434 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_39_44 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_39_446 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_39_449 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_39_468 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_39_471 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_39_483 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_39_491 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_39_497 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_39_50 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_39_503 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_39_505 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_39_509 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_39_512 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_39_53 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_39_534 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_39_537 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_39_551 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_39_554 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_39_561 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_39_610 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_39_613 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_39_623 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_39_626 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_39_638 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_39_642 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_39_645 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_39_65 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_39_650 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_39_653 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_39_656 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_39_659 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_39_662 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_39_665 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_39_668 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_39_671 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_39_673 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_39_676 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_39_679 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_39_68 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_39_713 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_39_80 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_39_95 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_39_98 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_3_108 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_3_169 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_3_288 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_3_3 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_3_31 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_3_315 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_3_322 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_3_328 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_3_332 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_3_337 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_3_343 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_3_355 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_3_367 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_3_379 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_3_391 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_3_393 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_3_405 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_3_415 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_3_418 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_3_421 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_3_430 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_3_537 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_3_558 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_3_57 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_3_609 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_3_66 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_3_713 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_3_86 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_3_91 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_40_111 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_40_124 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_40_133 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_40_136 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_40_141 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_40_149 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_40_154 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_40_166 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_40_178 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_40_190 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_40_193 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_40_200 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_40_203 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_40_215 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_40_227 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_40_232 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_40_251 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_40_256 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_40_259 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_40_294 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_40_3 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_40_306 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_40_309 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_40_317 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_40_322 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_40_329 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_40_341 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_40_388 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_40_391 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_40_394 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_40_406 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_40_418 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_40_421 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_40_431 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_40_434 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_40_445 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_40_457 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_40_461 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_40_464 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_40_475 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_40_477 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_40_524 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_40_533 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_40_536 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_40_54 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_40_542 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_40_562 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_40_580 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_40_583 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_40_586 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_40_598 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_40_631 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_40_634 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_40_638 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_40_641 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_40_650 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_40_658 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_40_66 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_40_677 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_40_699 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_40_75 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_40_78 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_40_81 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_40_93 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_40_96 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_40_99 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_41_101 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_41_109 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_41_136 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_41_140 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_41_15 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_41_164 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_41_167 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_41_169 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_41_191 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_41_209 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_41_212 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_41_225 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_41_229 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_41_253 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_41_265 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_41_275 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_41_278 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_41_281 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_41_3 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_41_304 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_41_337 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_41_349 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_41_353 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_41_385 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_41_393 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_41_396 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_41_399 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_41_40 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_41_426 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_41_429 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_41_432 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_41_446 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_41_449 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_41_46 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_41_461 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_41_466 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_41_472 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_41_475 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_41_502 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_41_513 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_41_525 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_41_537 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_41_54 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_41_554 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_41_557 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_41_561 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_41_57 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_41_575 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_41_578 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_41_581 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_41_585 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_41_594 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_41_597 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_41_603 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_41_625 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_41_629 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_41_632 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_41_655 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_41_713 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_41_86 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_41_89 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_42_101 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_42_104 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_42_123 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_42_126 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_42_138 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_42_141 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_42_145 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_42_15 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_42_173 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_42_176 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_42_190 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_42_193 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_42_213 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_42_225 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_42_233 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_42_251 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_42_253 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_42_256 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_42_268 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_42_27 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_42_272 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_42_29 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_42_290 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_42_293 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_42_3 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_42_305 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_42_32 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_42_340 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_42_344 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_42_347 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_42_358 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_42_393 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_42_424 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_42_427 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_42_43 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_42_448 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_42_451 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_42_454 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_42_466 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_42_47 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_42_470 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_42_473 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_42_477 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_42_50 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_42_511 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_42_523 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_42_531 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_42_533 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_42_537 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_42_544 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_42_547 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_42_559 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_42_562 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_42_568 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_42_571 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_42_575 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_42_578 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_42_581 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_42_584 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_42_587 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_42_594 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_42_597 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_42_600 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_42_603 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_42_61 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_42_610 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_42_613 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_42_616 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_42_622 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_42_625 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_42_628 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_42_631 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_42_643 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_42_65 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_42_68 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_42_699 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_42_74 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_42_93 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_43_111 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_43_125 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_43_137 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_43_149 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_43_15 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_43_156 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_43_165 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_43_169 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_43_181 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_43_213 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_43_216 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_43_225 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_43_254 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_43_257 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_43_260 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_43_268 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_43_27 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_43_278 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_43_284 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_43_287 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_43_290 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_43_3 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_43_304 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_43_325 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_43_328 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_43_337 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_43_343 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_43_346 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_43_35 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_43_357 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_43_360 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_43_364 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_43_378 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_43_381 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_43_384 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_43_387 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_43_393 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_43_40 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_43_422 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_43_426 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_43_429 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_43_434 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_43_437 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_43_449 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_43_45 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_43_465 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_43_468 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_43_474 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_43_477 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_43_480 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_43_484 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_43_492 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_43_495 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_43_503 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_43_505 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_43_517 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_43_526 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_43_529 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_43_53 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_43_532 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_43_535 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_43_547 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_43_555 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_43_559 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_43_566 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_43_569 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_43_57 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_43_573 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_43_576 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_43_579 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_43_582 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_43_586 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_43_589 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_43_592 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_43_595 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_43_598 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_43_601 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_43_604 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_43_615 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_43_622 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_43_625 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_43_628 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_43_631 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_43_634 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_43_637 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_43_640 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_43_645 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_43_648 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_43_69 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_43_705 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_43_77 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_43_96 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_43_99 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_44_100 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_44_135 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_44_139 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_44_141 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_44_15 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_44_166 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_44_178 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_44_192 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_44_195 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_44_206 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_44_218 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_44_226 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_44_253 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_44_265 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_44_27 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_44_290 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_44_294 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_44_297 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_44_3 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_44_309 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_44_312 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_44_322 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_44_334 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_44_346 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_44_358 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_44_365 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_44_377 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_44_381 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_44_392 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_44_417 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_44_421 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_44_427 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_44_435 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_44_439 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_44_449 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_44_452 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_44_464 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_44_468 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_44_477 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_44_489 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_44_497 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_44_500 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_44_514 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_44_517 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_44_52 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_44_528 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_44_531 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_44_533 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_44_536 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_44_539 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_44_542 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_44_546 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_44_549 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_44_553 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_44_559 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_44_562 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_44_565 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_44_568 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_44_573 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_44_576 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_44_579 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_44_582 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_44_585 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_44_589 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_44_592 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_44_604 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_44_625 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_44_632 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_44_635 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_44_638 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_44_64 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_44_641 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_44_645 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_44_648 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_44_71 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_44_74 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_44_85 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_44_88 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_45_106 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_45_113 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_45_124 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_45_127 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_45_139 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_45_147 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_45_15 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_45_159 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_45_163 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_45_166 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_45_169 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_45_181 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_45_203 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_45_215 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_45_22 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_45_223 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_45_225 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_45_244 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_45_247 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_45_259 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_45_26 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_45_278 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_45_281 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_45_289 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_45_29 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_45_294 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_45_297 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_45_3 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_45_308 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_45_317 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_45_329 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_45_335 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_45_337 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_45_349 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_45_35 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_45_361 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_45_373 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_45_391 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_45_393 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_45_396 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_45_399 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_45_402 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_45_405 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_45_408 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_45_420 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_45_432 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_45_444 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_45_449 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_45_461 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_45_471 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_45_479 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_45_482 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_45_485 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_45_491 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_45_494 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_45_500 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_45_503 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_45_505 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_45_508 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_45_511 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_45_515 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_45_518 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_45_521 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_45_525 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_45_528 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_45_53 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_45_531 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_45_534 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_45_553 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_45_556 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_45_559 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_45_561 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_45_566 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_45_569 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_45_57 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_45_574 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_45_577 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_45_580 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_45_587 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_45_590 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_45_595 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_45_598 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_45_603 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_45_606 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_45_609 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_45_612 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_45_615 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_45_617 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_45_620 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_45_623 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_45_628 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_45_631 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_45_713 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_45_91 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_45_94 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_46_100 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_46_103 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_46_107 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_46_110 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_46_121 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_46_124 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_46_136 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_46_141 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_46_145 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_46_164 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_46_176 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_46_188 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_46_195 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_46_205 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_46_208 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_46_211 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_46_214 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_46_238 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_46_241 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_46_251 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_46_253 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_46_265 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_46_269 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_46_272 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_46_284 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_46_296 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_46_3 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_46_309 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_46_332 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_46_344 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_46_356 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_46_365 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_46_377 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_46_38 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_46_394 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_46_397 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_46_408 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_46_411 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_46_419 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_46_421 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_46_433 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_46_439 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_46_442 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_46_445 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_46_456 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_46_459 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_46_462 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_46_465 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_46_468 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_46_471 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_46_477 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_46_480 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_46_490 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_46_50 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_46_514 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_46_517 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_46_520 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_46_528 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_46_531 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_46_533 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_46_536 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_46_539 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_46_542 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_46_555 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_46_560 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_46_567 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_46_570 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_46_573 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_46_62 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_46_626 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_46_645 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_46_83 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_46_93 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_46_97 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_47_107 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_47_110 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_47_113 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_47_118 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_47_123 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_47_135 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_47_141 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_47_144 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_47_164 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_47_167 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_47_169 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_47_181 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_47_205 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_47_208 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_47_216 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_47_221 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_47_228 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_47_246 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_47_249 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_47_292 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_47_3 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_47_304 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_47_312 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_47_337 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_47_349 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_47_361 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_47_369 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_47_381 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_47_384 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_47_393 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_47_397 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_47_400 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_47_439 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_47_442 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_47_449 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_47_453 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_47_456 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_47_46 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_47_467 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_47_472 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_47_475 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_47_49 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_47_508 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_47_511 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_47_522 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_47_533 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_47_545 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_47_548 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_47_55 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_47_551 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_47_554 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_47_557 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_47_561 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_47_564 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_47_567 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_47_57 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_47_570 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_47_605 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_47_61 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_47_670 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_47_68 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_47_71 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_48_108 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_48_133 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_48_139 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_48_141 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_48_15 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_48_173 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_48_181 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_48_189 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_48_193 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_48_214 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_48_222 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_48_234 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_48_238 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_48_250 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_48_253 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_48_259 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_48_26 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_48_262 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_48_288 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_48_3 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_48_300 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_48_309 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_48_312 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_48_340 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_48_343 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_48_355 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_48_37 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_48_388 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_48_40 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_48_405 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_48_408 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_48_411 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_48_419 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_48_421 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_48_429 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_48_432 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_48_443 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_48_446 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_48_449 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_48_452 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_48_455 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_48_470 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_48_473 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_48_477 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_48_48 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_48_51 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_48_513 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_48_567 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_48_585 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_48_610 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_48_63 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_48_677 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_48_710 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_48_75 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_48_83 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_49_111 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_49_116 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_49_135 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_49_140 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_49_15 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_49_151 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_49_163 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_49_166 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_49_169 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_49_208 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_49_211 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_49_214 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_49_225 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_49_235 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_49_239 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_49_242 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_49_248 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_49_279 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_49_289 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_49_292 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_49_296 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_49_3 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_49_334 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_49_337 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_49_340 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_49_352 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_49_360 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_49_365 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_49_377 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_49_380 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_49_40 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_49_414 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_49_422 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_49_425 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_49_447 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_49_457 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_49_460 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_49_463 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_49_466 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_49_469 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_49_472 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_49_475 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_49_495 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_49_498 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_49_501 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_49_505 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_49_55 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_49_556 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_49_559 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_49_569 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_49_57 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_49_588 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_49_591 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_49_670 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_49_68 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_49_72 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_49_75 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_49_81 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_49_84 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_4_104 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_4_107 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_4_154 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_4_307 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_4_319 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_4_327 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_4_340 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_4_352 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_4_365 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_4_377 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_4_38 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_4_389 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_4_401 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_4_413 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_4_419 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_4_421 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_4_424 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_4_430 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_4_500 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_4_530 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_4_549 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_4_587 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_4_592 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_4_642 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_4_713 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_4_78 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_4_85 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_50_110 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_50_127 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_50_130 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_50_134 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_50_137 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_50_141 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_50_145 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_50_15 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_50_151 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_50_154 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_50_166 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_50_178 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_50_182 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_50_194 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_50_205 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_50_208 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_50_216 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_50_243 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_50_246 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_50_253 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_50_256 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_50_27 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_50_276 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_50_279 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_50_29 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_50_291 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_50_299 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_50_3 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_50_302 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_50_305 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_50_317 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_50_334 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_50_360 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_50_363 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_50_365 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_50_397 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_50_400 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_50_41 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_50_415 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_50_421 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_50_429 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_50_432 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_50_454 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_50_457 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_50_460 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_50_470 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_50_493 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_50_496 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_50_508 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_50_511 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_50_520 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_50_529 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_50_533 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_50_536 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_50_578 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_50_589 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_50_643 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_50_65 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_50_661 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_50_699 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_50_713 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_50_77 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_50_83 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_50_85 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_51_113 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_51_116 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_51_121 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_51_124 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_51_136 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_51_161 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_51_167 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_51_169 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_51_181 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_51_189 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_51_194 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_51_206 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_51_218 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_51_225 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_51_245 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_51_248 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_51_260 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_51_264 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_51_273 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_51_279 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_51_281 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_51_293 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_51_3 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_51_307 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_51_335 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_51_34 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_51_354 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_51_357 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_51_373 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_51_378 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_51_381 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_51_384 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_51_387 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_51_391 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_51_393 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_51_405 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_51_408 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_51_411 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_51_414 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_51_417 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_51_445 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_51_449 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_51_46 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_51_502 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_51_54 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_51_558 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_51_609 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_51_670 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_51_713 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_51_74 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_51_86 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_51_94 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_52_115 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_52_118 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_52_121 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_52_124 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_52_136 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_52_141 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_52_15 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_52_162 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_52_165 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_52_173 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_52_178 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_52_181 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_52_19 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_52_192 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_52_195 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_52_197 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_52_209 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_52_233 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_52_242 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_52_246 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_52_249 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_52_253 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_52_265 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_52_277 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_52_289 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_52_3 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_52_301 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_52_307 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_52_309 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_52_32 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_52_331 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_52_337 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_52_349 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_52_36 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_52_361 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_52_365 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_52_373 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_52_377 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_52_389 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_52_397 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_52_401 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_52_404 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_52_407 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_52_417 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_52_48 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_52_525 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_52_586 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_52_60 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_52_642 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_52_66 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_52_698 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_52_701 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_52_704 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_52_713 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_52_78 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_52_85 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_52_97 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_53_100 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_53_108 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_53_113 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_53_117 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_53_120 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_53_123 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_53_131 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_53_136 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_53_139 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_53_15 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_53_158 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_53_161 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_53_167 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_53_169 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_53_181 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_53_187 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_53_191 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_53_194 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_53_197 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_53_202 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_53_206 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_53_209 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_53_212 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_53_225 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_53_228 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_53_23 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_53_234 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_53_239 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_53_242 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_53_245 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_53_248 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_53_251 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_53_254 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_53_257 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_53_262 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_53_274 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_53_281 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_53_293 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_53_299 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_53_3 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_53_303 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_53_306 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_53_309 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_53_312 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_53_315 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_53_326 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_53_329 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_53_332 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_53_337 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_53_34 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_53_347 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_53_359 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_53_362 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_53_365 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_53_368 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_53_371 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_53_374 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_53_386 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_53_398 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_53_401 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_53_405 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_53_45 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_53_48 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_53_503 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_53_558 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_53_57 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_53_615 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_53_670 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_53_685 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_53_69 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_53_73 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_53_76 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_53_88 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_54_130 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_54_133 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_54_137 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_54_141 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_54_144 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_54_147 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_54_15 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_54_152 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_54_155 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_54_158 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_54_166 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_54_169 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_54_173 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_54_177 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_54_192 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_54_208 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_54_21 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_54_211 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_54_215 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_54_219 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_54_222 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_54_225 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_54_230 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_54_233 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_54_236 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_54_239 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_54_25 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_54_251 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_54_256 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_54_259 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_54_264 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_54_267 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_54_270 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_54_277 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_54_281 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_54_29 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_54_297 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_54_3 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_54_302 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_54_305 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_54_328 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_54_332 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_54_341 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_54_361 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_54_365 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_54_370 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_54_373 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_54_376 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_54_379 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_54_382 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_54_387 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_54_390 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_54_41 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_54_410 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_54_474 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_54_493 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_54_53 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_54_586 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_54_643 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_54_661 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_54_69 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_54_698 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_54_713 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_54_73 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_54_76 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_54_80 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_54_83 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_54_85 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_54_89 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_55_11 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_55_122 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_55_155 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_55_158 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_55_162 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_55_165 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_55_169 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_55_214 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_55_223 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_55_3 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_55_304 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_55_308 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_55_311 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_55_335 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_55_35 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_55_38 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_55_385 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_55_446 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_55_50 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_55_528 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_55_53 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_55_547 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_55_551 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_55_614 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_55_633 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_55_671 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_55_678 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_55_80 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_55_83 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_55_86 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_56_15 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_56_172 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_56_21 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_56_25 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_56_251 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_56_253 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_56_3 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_56_307 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_56_326 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_56_350 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_56_46 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_56_474 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_56_530 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_56_586 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_56_642 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_56_698 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_56_85 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_56_88 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_56_91 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_56_94 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_57_11 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_57_110 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_57_148 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_57_213 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_57_222 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_57_225 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_57_243 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_57_252 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_57_278 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_57_290 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_57_3 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_57_302 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_57_334 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_57_337 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_57_446 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_57_449 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_57_452 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_57_47 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_57_50 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_57_501 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_57_53 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_57_558 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_57_561 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_57_613 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_57_670 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_57_673 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_57_676 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_57_91 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_57_96 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_57_99 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_58_149 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_58_15 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_58_164 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_58_19 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_58_197 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_58_211 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_58_227 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_58_231 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_58_247 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_58_251 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_58_278 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_58_283 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_58_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_58_3 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_58_44 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_58_474 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_58_530 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_58_586 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_58_642 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_58_698 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_58_710 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_58_83 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_58_91 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_59_11 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_59_113 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_59_141 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_59_160 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_59_207 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_59_253 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_59_275 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_59_279 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_59_281 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_59_3 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_59_309 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_59_337 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_59_341 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_59_369 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_59_391 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_59_419 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_59_447 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_59_449 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_59_452 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_59_474 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_59_502 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_59_505 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_59_508 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_59_530 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_59_558 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_59_561 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_59_564 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_59_57 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_59_586 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_59_614 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_59_617 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_59_620 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_59_642 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_59_670 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_59_673 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_59_698 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_59_713 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_5_102 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_5_140 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_5_225 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_5_241 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_5_278 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_5_293 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_5_312 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_5_318 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_5_330 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_5_337 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_5_349 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_5_361 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_5_373 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_5_385 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_5_391 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_5_393 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_5_405 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_5_417 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_5_423 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_5_426 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_5_429 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_5_446 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_5_449 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_5_46 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_5_68 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_5_713 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_6_11 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_6_227 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_6_251 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_6_268 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_6_285 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_6_288 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_6_29 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_6_307 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_6_312 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_6_324 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_6_33 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_6_336 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_6_348 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_6_360 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_6_365 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_6_377 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_6_389 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_6_401 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_6_406 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_6_418 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_6_421 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_6_425 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_6_475 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_6_493 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_6_530 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_6_536 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_6_585 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_6_713 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_6_96 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_6_99 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_7_102 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_7_119 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_7_201 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_7_223 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_7_256 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_7_266 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_7_295 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_7_306 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_7_312 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_7_333 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_7_337 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_7_349 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_7_353 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_7_359 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_7_371 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_7_383 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_7_387 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_7_390 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_7_424 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_7_432 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_7_465 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_7_468 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_7_471 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_7_505 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_7_508 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_7_511 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_7_556 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_7_612 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_7_642 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_7_645 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_7_648 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_7_666 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_7_73 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_7_76 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_8_130 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_8_179 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_8_223 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_8_234 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_8_261 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_8_273 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_8_281 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_8_295 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_8_3 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_8_307 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_8_309 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_8_317 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_8_338 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_8_350 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_8_362 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_8_365 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_8_381 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_8_384 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_8_387 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_8_405 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_8_417 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_8_432 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_8_459 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_8_470 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_8_473 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_8_480 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_8_58 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_8_61 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_8_621 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_8_643 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_8_653 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_8_701 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_8_713 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_8_75 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_9_113 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_9_169 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_9_214 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_9_270 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_9_3 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_9_300 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_9_334 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_9_340 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_9_343 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_9_351 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_9_355 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_9_358 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_9_381 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_9_391 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_9_401 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_9_404 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_9_407 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_9_428 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_9_436 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_9_447 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_9_549 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_9_593 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_9_620 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_9_649 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_9_713 ();
 sky130_fd_sc_hd__decap_3 PHY_0 ();
 sky130_fd_sc_hd__decap_3 PHY_1 ();
 sky130_fd_sc_hd__decap_3 PHY_10 ();
 sky130_fd_sc_hd__decap_3 PHY_100 ();
 sky130_fd_sc_hd__decap_3 PHY_101 ();
 sky130_fd_sc_hd__decap_3 PHY_102 ();
 sky130_fd_sc_hd__decap_3 PHY_103 ();
 sky130_fd_sc_hd__decap_3 PHY_104 ();
 sky130_fd_sc_hd__decap_3 PHY_105 ();
 sky130_fd_sc_hd__decap_3 PHY_106 ();
 sky130_fd_sc_hd__decap_3 PHY_107 ();
 sky130_fd_sc_hd__decap_3 PHY_108 ();
 sky130_fd_sc_hd__decap_3 PHY_109 ();
 sky130_fd_sc_hd__decap_3 PHY_11 ();
 sky130_fd_sc_hd__decap_3 PHY_110 ();
 sky130_fd_sc_hd__decap_3 PHY_111 ();
 sky130_fd_sc_hd__decap_3 PHY_112 ();
 sky130_fd_sc_hd__decap_3 PHY_113 ();
 sky130_fd_sc_hd__decap_3 PHY_114 ();
 sky130_fd_sc_hd__decap_3 PHY_115 ();
 sky130_fd_sc_hd__decap_3 PHY_116 ();
 sky130_fd_sc_hd__decap_3 PHY_117 ();
 sky130_fd_sc_hd__decap_3 PHY_118 ();
 sky130_fd_sc_hd__decap_3 PHY_119 ();
 sky130_fd_sc_hd__decap_3 PHY_12 ();
 sky130_fd_sc_hd__decap_3 PHY_13 ();
 sky130_fd_sc_hd__decap_3 PHY_14 ();
 sky130_fd_sc_hd__decap_3 PHY_15 ();
 sky130_fd_sc_hd__decap_3 PHY_16 ();
 sky130_fd_sc_hd__decap_3 PHY_17 ();
 sky130_fd_sc_hd__decap_3 PHY_18 ();
 sky130_fd_sc_hd__decap_3 PHY_19 ();
 sky130_fd_sc_hd__decap_3 PHY_2 ();
 sky130_fd_sc_hd__decap_3 PHY_20 ();
 sky130_fd_sc_hd__decap_3 PHY_21 ();
 sky130_fd_sc_hd__decap_3 PHY_22 ();
 sky130_fd_sc_hd__decap_3 PHY_23 ();
 sky130_fd_sc_hd__decap_3 PHY_24 ();
 sky130_fd_sc_hd__decap_3 PHY_25 ();
 sky130_fd_sc_hd__decap_3 PHY_26 ();
 sky130_fd_sc_hd__decap_3 PHY_27 ();
 sky130_fd_sc_hd__decap_3 PHY_28 ();
 sky130_fd_sc_hd__decap_3 PHY_29 ();
 sky130_fd_sc_hd__decap_3 PHY_3 ();
 sky130_fd_sc_hd__decap_3 PHY_30 ();
 sky130_fd_sc_hd__decap_3 PHY_31 ();
 sky130_fd_sc_hd__decap_3 PHY_32 ();
 sky130_fd_sc_hd__decap_3 PHY_33 ();
 sky130_fd_sc_hd__decap_3 PHY_34 ();
 sky130_fd_sc_hd__decap_3 PHY_35 ();
 sky130_fd_sc_hd__decap_3 PHY_36 ();
 sky130_fd_sc_hd__decap_3 PHY_37 ();
 sky130_fd_sc_hd__decap_3 PHY_38 ();
 sky130_fd_sc_hd__decap_3 PHY_39 ();
 sky130_fd_sc_hd__decap_3 PHY_4 ();
 sky130_fd_sc_hd__decap_3 PHY_40 ();
 sky130_fd_sc_hd__decap_3 PHY_41 ();
 sky130_fd_sc_hd__decap_3 PHY_42 ();
 sky130_fd_sc_hd__decap_3 PHY_43 ();
 sky130_fd_sc_hd__decap_3 PHY_44 ();
 sky130_fd_sc_hd__decap_3 PHY_45 ();
 sky130_fd_sc_hd__decap_3 PHY_46 ();
 sky130_fd_sc_hd__decap_3 PHY_47 ();
 sky130_fd_sc_hd__decap_3 PHY_48 ();
 sky130_fd_sc_hd__decap_3 PHY_49 ();
 sky130_fd_sc_hd__decap_3 PHY_5 ();
 sky130_fd_sc_hd__decap_3 PHY_50 ();
 sky130_fd_sc_hd__decap_3 PHY_51 ();
 sky130_fd_sc_hd__decap_3 PHY_52 ();
 sky130_fd_sc_hd__decap_3 PHY_53 ();
 sky130_fd_sc_hd__decap_3 PHY_54 ();
 sky130_fd_sc_hd__decap_3 PHY_55 ();
 sky130_fd_sc_hd__decap_3 PHY_56 ();
 sky130_fd_sc_hd__decap_3 PHY_57 ();
 sky130_fd_sc_hd__decap_3 PHY_58 ();
 sky130_fd_sc_hd__decap_3 PHY_59 ();
 sky130_fd_sc_hd__decap_3 PHY_6 ();
 sky130_fd_sc_hd__decap_3 PHY_60 ();
 sky130_fd_sc_hd__decap_3 PHY_61 ();
 sky130_fd_sc_hd__decap_3 PHY_62 ();
 sky130_fd_sc_hd__decap_3 PHY_63 ();
 sky130_fd_sc_hd__decap_3 PHY_64 ();
 sky130_fd_sc_hd__decap_3 PHY_65 ();
 sky130_fd_sc_hd__decap_3 PHY_66 ();
 sky130_fd_sc_hd__decap_3 PHY_67 ();
 sky130_fd_sc_hd__decap_3 PHY_68 ();
 sky130_fd_sc_hd__decap_3 PHY_69 ();
 sky130_fd_sc_hd__decap_3 PHY_7 ();
 sky130_fd_sc_hd__decap_3 PHY_70 ();
 sky130_fd_sc_hd__decap_3 PHY_71 ();
 sky130_fd_sc_hd__decap_3 PHY_72 ();
 sky130_fd_sc_hd__decap_3 PHY_73 ();
 sky130_fd_sc_hd__decap_3 PHY_74 ();
 sky130_fd_sc_hd__decap_3 PHY_75 ();
 sky130_fd_sc_hd__decap_3 PHY_76 ();
 sky130_fd_sc_hd__decap_3 PHY_77 ();
 sky130_fd_sc_hd__decap_3 PHY_78 ();
 sky130_fd_sc_hd__decap_3 PHY_79 ();
 sky130_fd_sc_hd__decap_3 PHY_8 ();
 sky130_fd_sc_hd__decap_3 PHY_80 ();
 sky130_fd_sc_hd__decap_3 PHY_81 ();
 sky130_fd_sc_hd__decap_3 PHY_82 ();
 sky130_fd_sc_hd__decap_3 PHY_83 ();
 sky130_fd_sc_hd__decap_3 PHY_84 ();
 sky130_fd_sc_hd__decap_3 PHY_85 ();
 sky130_fd_sc_hd__decap_3 PHY_86 ();
 sky130_fd_sc_hd__decap_3 PHY_87 ();
 sky130_fd_sc_hd__decap_3 PHY_88 ();
 sky130_fd_sc_hd__decap_3 PHY_89 ();
 sky130_fd_sc_hd__decap_3 PHY_9 ();
 sky130_fd_sc_hd__decap_3 PHY_90 ();
 sky130_fd_sc_hd__decap_3 PHY_91 ();
 sky130_fd_sc_hd__decap_3 PHY_92 ();
 sky130_fd_sc_hd__decap_3 PHY_93 ();
 sky130_fd_sc_hd__decap_3 PHY_94 ();
 sky130_fd_sc_hd__decap_3 PHY_95 ();
 sky130_fd_sc_hd__decap_3 PHY_96 ();
 sky130_fd_sc_hd__decap_3 PHY_97 ();
 sky130_fd_sc_hd__decap_3 PHY_98 ();
 sky130_fd_sc_hd__decap_3 PHY_99 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_120 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_121 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_122 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_123 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_124 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_125 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_126 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_127 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_128 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_129 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_130 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_131 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_132 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_133 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_134 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_135 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_136 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_137 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_138 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_139 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_140 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_141 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_142 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_143 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_144 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_145 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_146 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_147 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_148 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_149 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_150 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_151 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_152 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_153 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_154 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_155 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_156 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_157 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_158 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_159 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_160 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_161 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_162 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_163 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_164 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_165 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_166 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_167 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_168 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_169 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_170 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_171 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_172 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_173 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_174 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_175 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_176 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_177 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_178 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_179 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_180 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_181 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_182 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_183 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_184 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_185 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_186 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_187 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_188 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_189 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_190 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_191 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_192 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_193 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_194 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_195 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_196 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_197 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_198 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_199 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_200 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_201 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_202 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_203 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_204 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_205 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_206 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_207 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_208 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_209 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_210 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_211 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_212 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_213 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_214 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_215 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_216 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_217 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_218 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_219 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_220 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_221 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_222 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_223 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_224 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_225 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_226 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_227 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_228 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_229 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_230 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_231 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_232 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_233 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_234 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_235 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_236 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_237 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_238 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_239 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_240 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_241 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_242 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_243 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_244 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_245 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_246 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_247 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_248 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_249 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_250 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_251 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_252 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_253 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_254 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_255 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_256 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_257 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_258 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_259 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_260 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_261 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_262 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_263 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_264 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_265 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_266 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_267 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_268 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_269 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_270 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_271 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_272 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_273 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_274 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_275 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_276 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_277 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_278 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_279 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_280 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_281 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_282 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_283 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_284 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_285 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_286 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_287 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_288 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_289 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_290 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_291 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_292 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_293 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_294 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_295 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_296 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_297 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_298 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_299 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_300 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_301 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_302 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_303 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_304 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_305 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_306 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_307 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_308 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_309 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_310 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_311 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_312 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_313 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_314 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_315 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_316 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_317 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_318 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_319 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_320 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_321 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_322 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_323 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_324 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_325 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_326 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_327 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_328 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_329 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_330 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_331 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_332 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_333 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_334 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_335 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_336 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_337 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_338 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_339 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_340 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_341 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_342 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_343 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_344 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_345 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_346 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_347 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_348 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_349 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_350 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_351 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_352 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_353 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_354 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_355 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_356 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_357 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_358 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_359 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_360 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_361 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_362 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_363 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_364 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_365 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_366 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_367 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_368 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_369 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_370 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_371 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_372 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_373 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_374 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_375 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_376 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_377 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_378 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_379 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_380 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_381 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_382 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_383 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_384 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_385 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_386 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_387 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_388 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_389 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_390 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_391 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_392 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_393 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_394 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_395 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_396 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_397 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_398 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_399 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_400 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_401 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_402 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_403 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_404 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_405 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_406 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_407 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_408 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_409 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_410 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_411 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_412 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_413 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_414 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_415 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_416 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_417 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_418 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_419 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_420 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_421 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_422 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_423 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_424 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_425 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_426 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_427 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_428 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_429 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_430 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_431 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_432 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_433 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_434 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_435 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_436 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_437 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_438 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_439 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_440 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_441 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_442 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_443 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_444 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_445 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_446 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_447 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_448 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_449 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_450 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_451 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_452 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_453 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_454 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_455 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_456 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_457 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_458 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_459 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_460 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_461 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_462 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_463 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_464 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_465 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_466 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_467 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_468 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_469 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_470 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_471 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_472 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_473 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_474 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_475 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_476 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_477 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_478 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_479 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_480 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_481 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_482 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_483 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_484 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_485 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_486 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_487 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_488 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_489 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_490 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_491 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_492 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_493 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_494 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_495 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_496 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_497 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_498 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_499 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_500 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_501 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_502 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_503 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_504 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_505 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_506 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_507 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_508 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_509 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_510 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_511 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_512 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_513 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_514 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_515 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_516 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_517 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_518 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_519 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_520 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_521 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_522 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_523 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_524 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_525 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_526 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_527 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_528 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_529 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_530 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_531 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_532 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_533 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_534 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_535 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_536 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_537 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_538 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_539 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_540 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_541 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_542 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_543 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_544 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_545 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_546 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_547 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_548 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_549 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_550 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_551 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_552 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_553 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_554 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_555 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_556 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_557 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_558 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_559 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_560 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_561 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_562 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_563 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_564 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_565 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_566 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_567 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_568 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_569 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_570 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_571 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_572 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_573 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_574 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_575 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_576 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_577 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_578 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_579 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_580 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_581 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_582 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_583 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_584 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_585 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_586 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_587 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_588 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_589 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_590 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_591 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_592 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_593 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_594 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_595 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_596 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_597 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_598 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_599 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_600 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_601 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_602 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_603 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_604 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_605 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_606 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_607 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_608 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_609 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_610 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_611 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_612 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_613 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_614 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_615 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_616 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_617 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_618 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_619 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_620 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_621 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_622 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_623 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_624 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_625 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_626 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_627 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_628 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_629 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_630 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_631 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_632 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_633 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_634 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_635 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_636 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_637 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_638 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_639 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_640 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_641 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_642 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_643 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_644 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_645 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_646 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_647 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_648 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_649 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_650 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_651 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_652 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_653 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_654 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_655 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_656 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_657 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_658 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_659 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_660 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_661 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_662 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_663 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_664 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_665 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_666 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_667 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_668 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_669 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_670 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_671 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_672 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_673 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_674 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_675 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_676 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_677 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_678 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_679 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_680 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_681 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_682 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_683 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_684 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_685 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_686 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_687 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_688 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_689 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_690 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_691 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_692 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_693 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_694 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_695 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_696 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_697 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_698 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_699 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_700 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_701 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_702 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_703 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_704 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_705 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_706 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_707 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_708 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_709 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_710 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_711 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_712 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_713 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_714 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_715 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_716 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_717 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_718 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_719 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_720 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_721 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_722 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_723 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_724 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_725 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_726 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_727 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_728 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_729 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_730 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_731 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_732 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_733 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_734 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_735 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_736 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_737 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_738 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_739 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_740 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_741 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_742 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_743 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_744 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_745 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_746 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_747 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_748 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_749 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_750 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_751 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_752 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_753 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_754 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_755 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_756 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_757 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_758 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_759 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_760 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_761 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_762 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_763 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_764 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_765 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_766 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_767 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_768 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_769 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_770 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_771 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_772 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_773 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_774 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_775 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_776 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_777 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_778 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_779 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_780 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_781 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_782 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_783 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_784 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_785 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_786 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_787 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_788 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_789 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_790 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_791 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_792 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_793 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_794 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_795 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_796 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_797 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_798 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_799 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_800 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_801 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_802 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_803 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_804 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_805 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_806 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_807 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_808 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_809 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_810 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_811 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_812 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_813 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_814 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_815 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_816 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_817 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_818 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_819 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_820 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_821 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_822 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_823 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_824 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_825 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_826 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_827 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_828 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_829 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_830 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_831 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_832 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_833 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_834 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_835 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_836 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_837 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_838 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_839 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_840 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_841 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_842 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_843 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_844 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_845 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_846 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_847 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_848 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_849 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_850 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_851 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_852 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_853 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_854 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_855 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_856 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_857 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_858 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_859 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_860 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_861 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_862 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_863 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_864 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_865 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_866 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_867 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_868 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_869 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_870 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_871 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_872 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_873 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_874 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_875 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_876 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_877 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_878 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_879 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_880 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_881 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_882 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_883 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_884 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_885 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_886 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_887 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_888 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_889 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_890 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_891 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_892 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_893 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_894 ();
 sky130_fd_sc_hd__inv_2 _0952_ (.A(\current_state[1] ),
    .Y(_0004_));
 sky130_fd_sc_hd__inv_2 _0953_ (.A(net1209),
    .Y(_0520_));
 sky130_fd_sc_hd__inv_2 _0954_ (.A(net1167),
    .Y(_0521_));
 sky130_fd_sc_hd__inv_2 _0955_ (.A(updateRegs),
    .Y(_0522_));
 sky130_fd_sc_hd__inv_2 _0956_ (.A(net598),
    .Y(_0008_));
 sky130_fd_sc_hd__and2_2 _0957_ (.A(\current_state[0] ),
    .B(net591),
    .X(_0523_));
 sky130_fd_sc_hd__nand2_4 _0958_ (.A(\current_state[0] ),
    .B(net591),
    .Y(_0524_));
 sky130_fd_sc_hd__nor3_1 _0959_ (.A(net733),
    .B(net678),
    .C(net766),
    .Y(_0525_));
 sky130_fd_sc_hd__nor4_1 _0960_ (.A(net733),
    .B(net255),
    .C(net678),
    .D(net766),
    .Y(_0526_));
 sky130_fd_sc_hd__or4_2 _0961_ (.A(net733),
    .B(net255),
    .C(net678),
    .D(net766),
    .X(_0527_));
 sky130_fd_sc_hd__or2_2 _0962_ (.A(net1209),
    .B(net253),
    .X(_0528_));
 sky130_fd_sc_hd__or2_2 _0963_ (.A(_0527_),
    .B(_0528_),
    .X(_0529_));
 sky130_fd_sc_hd__or4_1 _0964_ (.A(net1142),
    .B(net1197),
    .C(net1084),
    .D(net1203),
    .X(_0530_));
 sky130_fd_sc_hd__or4b_1 _0965_ (.A(net1148),
    .B(net247),
    .C(net1216),
    .D_N(net692),
    .X(_0531_));
 sky130_fd_sc_hd__or4_2 _0966_ (.A(_0527_),
    .B(_0528_),
    .C(net1198),
    .D(net1217),
    .X(_0532_));
 sky130_fd_sc_hd__nand2_1 _0967_ (.A(net692),
    .B(net1148),
    .Y(_0533_));
 sky130_fd_sc_hd__or4_2 _0968_ (.A(net247),
    .B(_0527_),
    .C(_0528_),
    .D(net1149),
    .X(_0534_));
 sky130_fd_sc_hd__nor3_1 _0969_ (.A(net246),
    .B(net1198),
    .C(_0534_),
    .Y(_0535_));
 sky130_fd_sc_hd__and4b_1 _0970_ (.A_N(net247),
    .B(net246),
    .C(net692),
    .D(net1148),
    .X(_0536_));
 sky130_fd_sc_hd__or4b_1 _0971_ (.A(_0527_),
    .B(_0528_),
    .C(net1198),
    .D_N(_0536_),
    .X(_0537_));
 sky130_fd_sc_hd__or3_1 _0972_ (.A(net247),
    .B(net1216),
    .C(net1149),
    .X(_0538_));
 sky130_fd_sc_hd__or4_1 _0973_ (.A(net247),
    .B(_0529_),
    .C(_0530_),
    .D(net1149),
    .X(_0539_));
 sky130_fd_sc_hd__o211a_1 _0974_ (.A1(net1198),
    .A2(net1412),
    .B1(net1218),
    .C1(_0523_),
    .X(_0540_));
 sky130_fd_sc_hd__o211ai_1 _0975_ (.A1(net1198),
    .A2(_0534_),
    .B1(net1218),
    .C1(_0523_),
    .Y(_0541_));
 sky130_fd_sc_hd__and4_1 _0976_ (.A(net692),
    .B(net1148),
    .C(net247),
    .D(net1216),
    .X(_0542_));
 sky130_fd_sc_hd__nand4_1 _0977_ (.A(net692),
    .B(net1148),
    .C(net247),
    .D(net246),
    .Y(_0543_));
 sky130_fd_sc_hd__or3_1 _0978_ (.A(_0527_),
    .B(_0528_),
    .C(net693),
    .X(_0544_));
 sky130_fd_sc_hd__xor2_1 _0979_ (.A(net249),
    .B(net250),
    .X(_0545_));
 sky130_fd_sc_hd__or3b_1 _0980_ (.A(net1084),
    .B(_0545_),
    .C_N(net248),
    .X(_0546_));
 sky130_fd_sc_hd__or4bb_2 _0981_ (.A(net1084),
    .B(net1203),
    .C_N(net1142),
    .D_N(net1197),
    .X(_0547_));
 sky130_fd_sc_hd__nor2_1 _0982_ (.A(_0544_),
    .B(net1204),
    .Y(_0548_));
 sky130_fd_sc_hd__nor2_1 _0983_ (.A(net693),
    .B(_0547_),
    .Y(_0549_));
 sky130_fd_sc_hd__a311o_1 _0984_ (.A1(net1198),
    .A2(net1085),
    .A3(_0547_),
    .B1(net693),
    .C1(_0529_),
    .X(_0550_));
 sky130_fd_sc_hd__a311oi_1 _0985_ (.A1(net1198),
    .A2(net1085),
    .A3(_0547_),
    .B1(net693),
    .C1(_0529_),
    .Y(_0551_));
 sky130_fd_sc_hd__nor2_1 _0986_ (.A(net1199),
    .B(net1086),
    .Y(_0552_));
 sky130_fd_sc_hd__and4_1 _0987_ (.A(net1142),
    .B(net1197),
    .C(net1084),
    .D(net1203),
    .X(_0553_));
 sky130_fd_sc_hd__and2_2 _0988_ (.A(_0542_),
    .B(_0553_),
    .X(_0554_));
 sky130_fd_sc_hd__and2_1 _0989_ (.A(net1209),
    .B(net253),
    .X(_0555_));
 sky130_fd_sc_hd__and4_2 _0990_ (.A(_0526_),
    .B(_0542_),
    .C(_0553_),
    .D(net1439),
    .X(_0556_));
 sky130_fd_sc_hd__and3_1 _0991_ (.A(net1209),
    .B(net253),
    .C(net255),
    .X(_0557_));
 sky130_fd_sc_hd__and4_1 _0992_ (.A(net1209),
    .B(net253),
    .C(net733),
    .D(net255),
    .X(_0558_));
 sky130_fd_sc_hd__and4bb_1 _0993_ (.A_N(net678),
    .B_N(net766),
    .C(_0554_),
    .D(net1210),
    .X(_0559_));
 sky130_fd_sc_hd__o211a_1 _0994_ (.A1(net1440),
    .A2(net1211),
    .B1(_0540_),
    .C1(net694),
    .X(_0560_));
 sky130_fd_sc_hd__and4bb_2 _0995_ (.A_N(_0527_),
    .B_N(_0528_),
    .C(_0542_),
    .D(_0553_),
    .X(_0561_));
 sky130_fd_sc_hd__o21a_1 _0996_ (.A1(net1205),
    .A2(net1416),
    .B1(_0540_),
    .X(_0562_));
 sky130_fd_sc_hd__a32o_2 _0997_ (.A1(_0520_),
    .A2(net253),
    .A3(_0526_),
    .B1(_0557_),
    .B2(_0525_),
    .X(_0563_));
 sky130_fd_sc_hd__a211oi_4 _0998_ (.A1(_0554_),
    .A2(_0563_),
    .B1(_0561_),
    .C1(_0556_),
    .Y(_0564_));
 sky130_fd_sc_hd__and4b_1 _0999_ (.A_N(net678),
    .B(_0542_),
    .C(_0553_),
    .D(_0558_),
    .X(_0565_));
 sky130_fd_sc_hd__inv_2 _1000_ (.A(net679),
    .Y(_0566_));
 sky130_fd_sc_hd__o2bb2a_1 _1001_ (.A1_N(_0554_),
    .A2_N(_0563_),
    .B1(_0544_),
    .B2(net1085),
    .X(_0567_));
 sky130_fd_sc_hd__nand2_1 _1002_ (.A(net766),
    .B(net679),
    .Y(_0568_));
 sky130_fd_sc_hd__nor2_4 _1003_ (.A(\current_state[0] ),
    .B(net591),
    .Y(_0569_));
 sky130_fd_sc_hd__or2_2 _1004_ (.A(\current_state[0] ),
    .B(net591),
    .X(_0570_));
 sky130_fd_sc_hd__and4bb_1 _1005_ (.A_N(net879),
    .B_N(net932),
    .C(net900),
    .D(net946),
    .X(_0571_));
 sky130_fd_sc_hd__and4b_1 _1006_ (.A_N(net904),
    .B(net893),
    .C(net864),
    .D(net783),
    .X(_0572_));
 sky130_fd_sc_hd__nand2_2 _1007_ (.A(_0571_),
    .B(_0572_),
    .Y(_0573_));
 sky130_fd_sc_hd__nand2_1 _1008_ (.A(net560),
    .B(_0573_),
    .Y(_0574_));
 sky130_fd_sc_hd__a21o_1 _1009_ (.A1(net1218),
    .A2(_0537_),
    .B1(_0524_),
    .X(_0575_));
 sky130_fd_sc_hd__o211ai_1 _1010_ (.A1(net1199),
    .A2(_0567_),
    .B1(_0574_),
    .C1(_0575_),
    .Y(_0576_));
 sky130_fd_sc_hd__and2b_1 _1011_ (.A_N(net766),
    .B(net678),
    .X(_0577_));
 sky130_fd_sc_hd__and4b_1 _1012_ (.A_N(_0577_),
    .B(_0558_),
    .C(_0553_),
    .D(_0542_),
    .X(_0578_));
 sky130_fd_sc_hd__a2111o_1 _1013_ (.A1(_0554_),
    .A2(_0563_),
    .B1(_0578_),
    .C1(_0556_),
    .D1(_0561_),
    .X(_0579_));
 sky130_fd_sc_hd__nand4_1 _1014_ (.A(net733),
    .B(net255),
    .C(_0554_),
    .D(_0555_),
    .Y(_0580_));
 sky130_fd_sc_hd__o21a_1 _1015_ (.A1(_0577_),
    .A2(net734),
    .B1(_0564_),
    .X(_0581_));
 sky130_fd_sc_hd__a211o_1 _1016_ (.A1(net767),
    .A2(_0579_),
    .B1(net1199),
    .C1(net1086),
    .X(_0582_));
 sky130_fd_sc_hd__o21ba_1 _1017_ (.A1(_0549_),
    .A2(_0554_),
    .B1_N(_0529_),
    .X(_0583_));
 sky130_fd_sc_hd__a211oi_1 _1018_ (.A1(_0538_),
    .A2(net693),
    .B1(_0529_),
    .C1(net1198),
    .Y(_0584_));
 sky130_fd_sc_hd__a32o_1 _1019_ (.A1(_0523_),
    .A2(net1218),
    .A3(net1435),
    .B1(_0583_),
    .B2(_0540_),
    .X(_0585_));
 sky130_fd_sc_hd__o2111a_1 _1020_ (.A1(net678),
    .A2(net734),
    .B1(_0564_),
    .C1(net694),
    .D1(net1150),
    .X(_0586_));
 sky130_fd_sc_hd__or4b_1 _1021_ (.A(net695),
    .B(_0576_),
    .C(net1219),
    .D_N(net1087),
    .X(_0587_));
 sky130_fd_sc_hd__or2_1 _1022_ (.A(net595),
    .B(net1088),
    .X(_0588_));
 sky130_fd_sc_hd__nor2_2 _1023_ (.A(_0570_),
    .B(_0573_),
    .Y(_0589_));
 sky130_fd_sc_hd__nor4_1 _1024_ (.A(net1177),
    .B(net1185),
    .C(net1192),
    .D(net1181),
    .Y(_0590_));
 sky130_fd_sc_hd__nor2_1 _1025_ (.A(net777),
    .B(net1167),
    .Y(_0591_));
 sky130_fd_sc_hd__and3_4 _1026_ (.A(net745),
    .B(_0590_),
    .C(net778),
    .X(_0592_));
 sky130_fd_sc_hd__nand3_1 _1027_ (.A(net745),
    .B(_0590_),
    .C(net778),
    .Y(_0593_));
 sky130_fd_sc_hd__mux2_1 _1028_ (.A0(\reg_temp[162] ),
    .A1(net1447),
    .S(net590),
    .X(_0594_));
 sky130_fd_sc_hd__a22o_1 _1029_ (.A1(net1240),
    .A2(net532),
    .B1(net557),
    .B2(net1448),
    .X(_0519_));
 sky130_fd_sc_hd__mux2_1 _1030_ (.A0(\reg_temp[161] ),
    .A1(net1445),
    .S(net590),
    .X(_0595_));
 sky130_fd_sc_hd__a22o_1 _1031_ (.A1(net1245),
    .A2(net532),
    .B1(net557),
    .B2(net1446),
    .X(_0518_));
 sky130_fd_sc_hd__mux2_1 _1032_ (.A0(\reg_temp[160] ),
    .A1(\reg_temp[78] ),
    .S(net590),
    .X(_0596_));
 sky130_fd_sc_hd__a22o_1 _1033_ (.A1(net1244),
    .A2(net532),
    .B1(net557),
    .B2(_0596_),
    .X(_0517_));
 sky130_fd_sc_hd__mux2_1 _1034_ (.A0(\reg_temp[159] ),
    .A1(\reg_temp[77] ),
    .S(net590),
    .X(_0597_));
 sky130_fd_sc_hd__a22o_1 _1035_ (.A1(net1256),
    .A2(net532),
    .B1(net556),
    .B2(_0597_),
    .X(_0516_));
 sky130_fd_sc_hd__mux2_1 _1036_ (.A0(\reg_temp[158] ),
    .A1(\reg_temp[76] ),
    .S(net589),
    .X(_0598_));
 sky130_fd_sc_hd__a22o_1 _1037_ (.A1(net1294),
    .A2(net531),
    .B1(net556),
    .B2(_0598_),
    .X(_0515_));
 sky130_fd_sc_hd__mux2_2 _1038_ (.A0(\reg_temp[157] ),
    .A1(\reg_temp[75] ),
    .S(_0592_),
    .X(_0599_));
 sky130_fd_sc_hd__a22o_1 _1039_ (.A1(net1228),
    .A2(net532),
    .B1(net557),
    .B2(_0599_),
    .X(_0514_));
 sky130_fd_sc_hd__mux2_1 _1040_ (.A0(\reg_temp[156] ),
    .A1(\reg_temp[74] ),
    .S(net590),
    .X(_0600_));
 sky130_fd_sc_hd__a22o_1 _1041_ (.A1(net1259),
    .A2(net532),
    .B1(net557),
    .B2(_0600_),
    .X(_0513_));
 sky130_fd_sc_hd__mux2_1 _1042_ (.A0(\reg_temp[155] ),
    .A1(\reg_temp[73] ),
    .S(net590),
    .X(_0601_));
 sky130_fd_sc_hd__a22o_1 _1043_ (.A1(net1253),
    .A2(net532),
    .B1(net557),
    .B2(_0601_),
    .X(_0512_));
 sky130_fd_sc_hd__mux2_1 _1044_ (.A0(\reg_temp[154] ),
    .A1(\reg_temp[72] ),
    .S(net589),
    .X(_0602_));
 sky130_fd_sc_hd__a22o_1 _1045_ (.A1(net1307),
    .A2(net531),
    .B1(net556),
    .B2(_0602_),
    .X(_0511_));
 sky130_fd_sc_hd__mux2_1 _1046_ (.A0(\reg_temp[153] ),
    .A1(\reg_temp[71] ),
    .S(net590),
    .X(_0603_));
 sky130_fd_sc_hd__a22o_1 _1047_ (.A1(net1252),
    .A2(net532),
    .B1(net557),
    .B2(_0603_),
    .X(_0510_));
 sky130_fd_sc_hd__mux2_1 _1048_ (.A0(\reg_temp[152] ),
    .A1(\reg_temp[70] ),
    .S(net590),
    .X(_0604_));
 sky130_fd_sc_hd__a22o_1 _1049_ (.A1(net1251),
    .A2(net531),
    .B1(net556),
    .B2(_0604_),
    .X(_0509_));
 sky130_fd_sc_hd__mux2_1 _1050_ (.A0(\reg_temp[151] ),
    .A1(\reg_temp[69] ),
    .S(net590),
    .X(_0605_));
 sky130_fd_sc_hd__a22o_1 _1051_ (.A1(net1249),
    .A2(net532),
    .B1(net557),
    .B2(_0605_),
    .X(_0508_));
 sky130_fd_sc_hd__mux2_1 _1052_ (.A0(\reg_temp[150] ),
    .A1(\reg_temp[68] ),
    .S(net590),
    .X(_0606_));
 sky130_fd_sc_hd__a22o_1 _1053_ (.A1(net1248),
    .A2(net532),
    .B1(net557),
    .B2(_0606_),
    .X(_0507_));
 sky130_fd_sc_hd__mux2_1 _1054_ (.A0(\reg_temp[149] ),
    .A1(\reg_temp[67] ),
    .S(net590),
    .X(_0607_));
 sky130_fd_sc_hd__a22o_1 _1055_ (.A1(net1247),
    .A2(net531),
    .B1(net557),
    .B2(_0607_),
    .X(_0506_));
 sky130_fd_sc_hd__mux2_1 _1056_ (.A0(\reg_temp[148] ),
    .A1(\reg_temp[66] ),
    .S(net590),
    .X(_0608_));
 sky130_fd_sc_hd__a22o_1 _1057_ (.A1(net1246),
    .A2(net532),
    .B1(net557),
    .B2(_0608_),
    .X(_0505_));
 sky130_fd_sc_hd__mux2_1 _1058_ (.A0(\reg_temp[147] ),
    .A1(\reg_temp[65] ),
    .S(net590),
    .X(_0609_));
 sky130_fd_sc_hd__a22o_1 _1059_ (.A1(net1230),
    .A2(net533),
    .B1(net558),
    .B2(_0609_),
    .X(_0504_));
 sky130_fd_sc_hd__mux2_1 _1060_ (.A0(\reg_temp[146] ),
    .A1(\reg_temp[64] ),
    .S(net589),
    .X(_0610_));
 sky130_fd_sc_hd__a22o_1 _1061_ (.A1(net1301),
    .A2(net531),
    .B1(net556),
    .B2(_0610_),
    .X(_0503_));
 sky130_fd_sc_hd__mux2_1 _1062_ (.A0(\reg_temp[145] ),
    .A1(\reg_temp[63] ),
    .S(net589),
    .X(_0611_));
 sky130_fd_sc_hd__a22o_1 _1063_ (.A1(net1235),
    .A2(net533),
    .B1(net558),
    .B2(_0611_),
    .X(_0502_));
 sky130_fd_sc_hd__mux2_1 _1064_ (.A0(\reg_temp[144] ),
    .A1(\reg_temp[62] ),
    .S(net589),
    .X(_0612_));
 sky130_fd_sc_hd__a22o_1 _1065_ (.A1(net1308),
    .A2(net531),
    .B1(net556),
    .B2(_0612_),
    .X(_0501_));
 sky130_fd_sc_hd__mux2_1 _1066_ (.A0(\reg_temp[143] ),
    .A1(\reg_temp[61] ),
    .S(net589),
    .X(_0613_));
 sky130_fd_sc_hd__a22o_1 _1067_ (.A1(net508),
    .A2(net531),
    .B1(net556),
    .B2(_0613_),
    .X(_0500_));
 sky130_fd_sc_hd__mux2_1 _1068_ (.A0(\reg_temp[142] ),
    .A1(\reg_temp[60] ),
    .S(net589),
    .X(_0614_));
 sky130_fd_sc_hd__a22o_1 _1069_ (.A1(net1233),
    .A2(net533),
    .B1(net558),
    .B2(_0614_),
    .X(_0499_));
 sky130_fd_sc_hd__mux2_1 _1070_ (.A0(\reg_temp[141] ),
    .A1(\reg_temp[59] ),
    .S(net589),
    .X(_0615_));
 sky130_fd_sc_hd__a22o_1 _1071_ (.A1(net1232),
    .A2(net533),
    .B1(net558),
    .B2(_0615_),
    .X(_0498_));
 sky130_fd_sc_hd__mux2_1 _1072_ (.A0(\reg_temp[140] ),
    .A1(net1651),
    .S(net589),
    .X(_0616_));
 sky130_fd_sc_hd__a22o_1 _1073_ (.A1(net1302),
    .A2(net531),
    .B1(net556),
    .B2(_0616_),
    .X(_0497_));
 sky130_fd_sc_hd__mux2_1 _1074_ (.A0(\reg_temp[139] ),
    .A1(\reg_temp[57] ),
    .S(net589),
    .X(_0617_));
 sky130_fd_sc_hd__a22o_1 _1075_ (.A1(net1293),
    .A2(net531),
    .B1(net556),
    .B2(_0617_),
    .X(_0496_));
 sky130_fd_sc_hd__mux2_2 _1076_ (.A0(\reg_temp[138] ),
    .A1(\reg_temp[56] ),
    .S(net589),
    .X(_0618_));
 sky130_fd_sc_hd__a22o_1 _1077_ (.A1(net1289),
    .A2(net531),
    .B1(net556),
    .B2(_0618_),
    .X(_0495_));
 sky130_fd_sc_hd__mux2_1 _1078_ (.A0(\reg_temp[137] ),
    .A1(\reg_temp[55] ),
    .S(net589),
    .X(_0619_));
 sky130_fd_sc_hd__a22o_1 _1079_ (.A1(net1292),
    .A2(net531),
    .B1(net556),
    .B2(_0619_),
    .X(_0494_));
 sky130_fd_sc_hd__mux2_1 _1080_ (.A0(\reg_temp[136] ),
    .A1(\reg_temp[54] ),
    .S(net589),
    .X(_0620_));
 sky130_fd_sc_hd__a22o_1 _1081_ (.A1(net501),
    .A2(net531),
    .B1(net556),
    .B2(_0620_),
    .X(_0493_));
 sky130_fd_sc_hd__mux2_1 _1082_ (.A0(\reg_temp[135] ),
    .A1(\reg_temp[53] ),
    .S(net589),
    .X(_0621_));
 sky130_fd_sc_hd__a22o_1 _1083_ (.A1(net500),
    .A2(net531),
    .B1(net556),
    .B2(_0621_),
    .X(_0492_));
 sky130_fd_sc_hd__mux2_1 _1084_ (.A0(\reg_temp[134] ),
    .A1(\reg_temp[52] ),
    .S(net589),
    .X(_0622_));
 sky130_fd_sc_hd__a22o_1 _1085_ (.A1(net1309),
    .A2(net531),
    .B1(net556),
    .B2(_0622_),
    .X(_0491_));
 sky130_fd_sc_hd__mux2_1 _1086_ (.A0(\reg_temp[133] ),
    .A1(\reg_temp[51] ),
    .S(net589),
    .X(_0623_));
 sky130_fd_sc_hd__a22o_1 _1087_ (.A1(net498),
    .A2(net531),
    .B1(net556),
    .B2(_0623_),
    .X(_0490_));
 sky130_fd_sc_hd__mux2_1 _1088_ (.A0(\reg_temp[132] ),
    .A1(\reg_temp[50] ),
    .S(net588),
    .X(_0624_));
 sky130_fd_sc_hd__a22o_1 _1089_ (.A1(net1237),
    .A2(net533),
    .B1(net558),
    .B2(_0624_),
    .X(_0489_));
 sky130_fd_sc_hd__mux2_1 _1090_ (.A0(net1444),
    .A1(\reg_temp[49] ),
    .S(net590),
    .X(_0625_));
 sky130_fd_sc_hd__a22o_1 _1091_ (.A1(net1231),
    .A2(net533),
    .B1(net558),
    .B2(_0625_),
    .X(_0488_));
 sky130_fd_sc_hd__mux2_1 _1092_ (.A0(\reg_temp[130] ),
    .A1(\reg_temp[48] ),
    .S(net585),
    .X(_0626_));
 sky130_fd_sc_hd__a22o_1 _1093_ (.A1(net1236),
    .A2(net533),
    .B1(net558),
    .B2(_0626_),
    .X(_0487_));
 sky130_fd_sc_hd__mux2_1 _1094_ (.A0(\reg_temp[129] ),
    .A1(\reg_temp[47] ),
    .S(net590),
    .X(_0627_));
 sky130_fd_sc_hd__a22o_1 _1095_ (.A1(net1243),
    .A2(net531),
    .B1(net556),
    .B2(_0627_),
    .X(_0486_));
 sky130_fd_sc_hd__mux2_1 _1096_ (.A0(\reg_temp[128] ),
    .A1(net1449),
    .S(net588),
    .X(_0628_));
 sky130_fd_sc_hd__a22o_1 _1097_ (.A1(net1229),
    .A2(net533),
    .B1(net558),
    .B2(_0628_),
    .X(_0485_));
 sky130_fd_sc_hd__mux2_1 _1098_ (.A0(\reg_temp[127] ),
    .A1(\reg_temp[45] ),
    .S(net588),
    .X(_0629_));
 sky130_fd_sc_hd__a22o_1 _1099_ (.A1(net1223),
    .A2(net530),
    .B1(net555),
    .B2(_0629_),
    .X(_0484_));
 sky130_fd_sc_hd__mux2_1 _1100_ (.A0(\reg_temp[126] ),
    .A1(\reg_temp[44] ),
    .S(net585),
    .X(_0630_));
 sky130_fd_sc_hd__a22o_1 _1101_ (.A1(net491),
    .A2(net528),
    .B1(net553),
    .B2(_0630_),
    .X(_0483_));
 sky130_fd_sc_hd__mux2_1 _1102_ (.A0(\reg_temp[125] ),
    .A1(\reg_temp[43] ),
    .S(net588),
    .X(_0631_));
 sky130_fd_sc_hd__a22o_1 _1103_ (.A1(net1250),
    .A2(net528),
    .B1(net553),
    .B2(_0631_),
    .X(_0482_));
 sky130_fd_sc_hd__mux2_1 _1104_ (.A0(\reg_temp[124] ),
    .A1(\reg_temp[42] ),
    .S(net585),
    .X(_0632_));
 sky130_fd_sc_hd__a22o_1 _1105_ (.A1(net1277),
    .A2(net528),
    .B1(net553),
    .B2(_0632_),
    .X(_0481_));
 sky130_fd_sc_hd__mux2_1 _1106_ (.A0(net1633),
    .A1(\reg_temp[41] ),
    .S(net585),
    .X(_0633_));
 sky130_fd_sc_hd__a22o_1 _1107_ (.A1(net1420),
    .A2(net528),
    .B1(net553),
    .B2(_0633_),
    .X(_0480_));
 sky130_fd_sc_hd__mux2_1 _1108_ (.A0(\reg_temp[122] ),
    .A1(\reg_temp[40] ),
    .S(net585),
    .X(_0634_));
 sky130_fd_sc_hd__a22o_1 _1109_ (.A1(net487),
    .A2(net528),
    .B1(net553),
    .B2(_0634_),
    .X(_0479_));
 sky130_fd_sc_hd__mux2_1 _1110_ (.A0(\reg_temp[121] ),
    .A1(\reg_temp[39] ),
    .S(net588),
    .X(_0635_));
 sky130_fd_sc_hd__a22o_1 _1111_ (.A1(net1242),
    .A2(net528),
    .B1(net553),
    .B2(_0635_),
    .X(_0478_));
 sky130_fd_sc_hd__mux2_1 _1112_ (.A0(\reg_temp[120] ),
    .A1(\reg_temp[38] ),
    .S(net588),
    .X(_0636_));
 sky130_fd_sc_hd__a22o_1 _1113_ (.A1(net1241),
    .A2(net529),
    .B1(net554),
    .B2(_0636_),
    .X(_0477_));
 sky130_fd_sc_hd__mux2_1 _1114_ (.A0(\reg_temp[119] ),
    .A1(\reg_temp[37] ),
    .S(net586),
    .X(_0637_));
 sky130_fd_sc_hd__a22o_1 _1115_ (.A1(net1303),
    .A2(net529),
    .B1(net554),
    .B2(_0637_),
    .X(_0476_));
 sky130_fd_sc_hd__mux2_1 _1116_ (.A0(\reg_temp[118] ),
    .A1(\reg_temp[36] ),
    .S(net586),
    .X(_0638_));
 sky130_fd_sc_hd__a22o_1 _1117_ (.A1(net1306),
    .A2(net529),
    .B1(net554),
    .B2(_0638_),
    .X(_0475_));
 sky130_fd_sc_hd__mux2_1 _1118_ (.A0(\reg_temp[117] ),
    .A1(\reg_temp[35] ),
    .S(net587),
    .X(_0639_));
 sky130_fd_sc_hd__a22o_1 _1119_ (.A1(net1305),
    .A2(net527),
    .B1(net552),
    .B2(_0639_),
    .X(_0474_));
 sky130_fd_sc_hd__mux2_1 _1120_ (.A0(\reg_temp[116] ),
    .A1(\reg_temp[34] ),
    .S(net586),
    .X(_0640_));
 sky130_fd_sc_hd__a22o_1 _1121_ (.A1(net1300),
    .A2(net527),
    .B1(net552),
    .B2(_0640_),
    .X(_0473_));
 sky130_fd_sc_hd__mux2_1 _1122_ (.A0(\reg_temp[115] ),
    .A1(\reg_temp[33] ),
    .S(net586),
    .X(_0641_));
 sky130_fd_sc_hd__a22o_1 _1123_ (.A1(net1304),
    .A2(net529),
    .B1(net554),
    .B2(_0641_),
    .X(_0472_));
 sky130_fd_sc_hd__mux2_1 _1124_ (.A0(\reg_temp[114] ),
    .A1(\reg_temp[32] ),
    .S(net587),
    .X(_0642_));
 sky130_fd_sc_hd__a22o_1 _1125_ (.A1(net1299),
    .A2(net529),
    .B1(net554),
    .B2(_0642_),
    .X(_0471_));
 sky130_fd_sc_hd__mux2_1 _1126_ (.A0(\reg_temp[113] ),
    .A1(\reg_temp[31] ),
    .S(net587),
    .X(_0643_));
 sky130_fd_sc_hd__a22o_1 _1127_ (.A1(net1272),
    .A2(net527),
    .B1(net552),
    .B2(_0643_),
    .X(_0470_));
 sky130_fd_sc_hd__mux2_1 _1128_ (.A0(\reg_temp[112] ),
    .A1(\reg_temp[30] ),
    .S(net587),
    .X(_0644_));
 sky130_fd_sc_hd__a22o_1 _1129_ (.A1(net477),
    .A2(net527),
    .B1(net552),
    .B2(_0644_),
    .X(_0469_));
 sky130_fd_sc_hd__mux2_1 _1130_ (.A0(\reg_temp[111] ),
    .A1(\reg_temp[29] ),
    .S(net587),
    .X(_0645_));
 sky130_fd_sc_hd__a22o_1 _1131_ (.A1(net1255),
    .A2(net528),
    .B1(net553),
    .B2(_0645_),
    .X(_0468_));
 sky130_fd_sc_hd__mux2_1 _1132_ (.A0(\reg_temp[110] ),
    .A1(\reg_temp[28] ),
    .S(net587),
    .X(_0646_));
 sky130_fd_sc_hd__a22o_1 _1133_ (.A1(net475),
    .A2(net529),
    .B1(net555),
    .B2(_0646_),
    .X(_0467_));
 sky130_fd_sc_hd__mux2_1 _1134_ (.A0(\reg_temp[109] ),
    .A1(\reg_temp[27] ),
    .S(net587),
    .X(_0647_));
 sky130_fd_sc_hd__a22o_1 _1135_ (.A1(net1271),
    .A2(net530),
    .B1(net554),
    .B2(_0647_),
    .X(_0466_));
 sky130_fd_sc_hd__mux2_1 _1136_ (.A0(\reg_temp[108] ),
    .A1(\reg_temp[26] ),
    .S(net587),
    .X(_0648_));
 sky130_fd_sc_hd__a22o_1 _1137_ (.A1(net473),
    .A2(net528),
    .B1(net553),
    .B2(_0648_),
    .X(_0465_));
 sky130_fd_sc_hd__mux2_1 _1138_ (.A0(\reg_temp[107] ),
    .A1(\reg_temp[25] ),
    .S(net587),
    .X(_0649_));
 sky130_fd_sc_hd__a22o_1 _1139_ (.A1(net1254),
    .A2(net528),
    .B1(net553),
    .B2(_0649_),
    .X(_0464_));
 sky130_fd_sc_hd__mux2_1 _1140_ (.A0(\reg_temp[106] ),
    .A1(\reg_temp[24] ),
    .S(net586),
    .X(_0650_));
 sky130_fd_sc_hd__a22o_1 _1141_ (.A1(net471),
    .A2(net527),
    .B1(net552),
    .B2(_0650_),
    .X(_0463_));
 sky130_fd_sc_hd__mux2_1 _1142_ (.A0(\reg_temp[105] ),
    .A1(\reg_temp[23] ),
    .S(net586),
    .X(_0651_));
 sky130_fd_sc_hd__a22o_1 _1143_ (.A1(net1273),
    .A2(net527),
    .B1(net552),
    .B2(_0651_),
    .X(_0462_));
 sky130_fd_sc_hd__mux2_1 _1144_ (.A0(\reg_temp[104] ),
    .A1(\reg_temp[22] ),
    .S(net587),
    .X(_0652_));
 sky130_fd_sc_hd__a22o_1 _1145_ (.A1(net469),
    .A2(net530),
    .B1(net555),
    .B2(_0652_),
    .X(_0461_));
 sky130_fd_sc_hd__mux2_1 _1146_ (.A0(\reg_temp[103] ),
    .A1(\reg_temp[21] ),
    .S(net586),
    .X(_0653_));
 sky130_fd_sc_hd__a22o_1 _1147_ (.A1(net1274),
    .A2(net527),
    .B1(net552),
    .B2(_0653_),
    .X(_0460_));
 sky130_fd_sc_hd__mux2_1 _1148_ (.A0(\reg_temp[102] ),
    .A1(\reg_temp[20] ),
    .S(net586),
    .X(_0654_));
 sky130_fd_sc_hd__a22o_1 _1149_ (.A1(net1296),
    .A2(net529),
    .B1(net554),
    .B2(_0654_),
    .X(_0459_));
 sky130_fd_sc_hd__mux2_1 _1150_ (.A0(\reg_temp[101] ),
    .A1(\reg_temp[19] ),
    .S(net586),
    .X(_0655_));
 sky130_fd_sc_hd__a22o_1 _1151_ (.A1(net1283),
    .A2(net529),
    .B1(net554),
    .B2(_0655_),
    .X(_0458_));
 sky130_fd_sc_hd__mux2_1 _1152_ (.A0(\reg_temp[100] ),
    .A1(\reg_temp[18] ),
    .S(net586),
    .X(_0656_));
 sky130_fd_sc_hd__a22o_1 _1153_ (.A1(net1227),
    .A2(net530),
    .B1(net555),
    .B2(_0656_),
    .X(_0457_));
 sky130_fd_sc_hd__mux2_1 _1154_ (.A0(\reg_temp[99] ),
    .A1(\reg_temp[17] ),
    .S(net586),
    .X(_0657_));
 sky130_fd_sc_hd__a22o_1 _1155_ (.A1(net1264),
    .A2(net527),
    .B1(net552),
    .B2(_0657_),
    .X(_0456_));
 sky130_fd_sc_hd__mux2_1 _1156_ (.A0(\reg_temp[98] ),
    .A1(\reg_temp[16] ),
    .S(net587),
    .X(_0658_));
 sky130_fd_sc_hd__a22o_1 _1157_ (.A1(net1224),
    .A2(net530),
    .B1(net555),
    .B2(_0658_),
    .X(_0455_));
 sky130_fd_sc_hd__mux2_1 _1158_ (.A0(\reg_temp[97] ),
    .A1(\reg_temp[15] ),
    .S(net586),
    .X(_0659_));
 sky130_fd_sc_hd__a22o_1 _1159_ (.A1(net1263),
    .A2(net527),
    .B1(net552),
    .B2(_0659_),
    .X(_0454_));
 sky130_fd_sc_hd__mux2_1 _1160_ (.A0(\reg_temp[96] ),
    .A1(\reg_temp[14] ),
    .S(net586),
    .X(_0660_));
 sky130_fd_sc_hd__a22o_1 _1161_ (.A1(net461),
    .A2(net527),
    .B1(net552),
    .B2(_0660_),
    .X(_0453_));
 sky130_fd_sc_hd__mux2_1 _1162_ (.A0(\reg_temp[95] ),
    .A1(\reg_temp[13] ),
    .S(net585),
    .X(_0661_));
 sky130_fd_sc_hd__a22o_1 _1163_ (.A1(net1297),
    .A2(net529),
    .B1(net554),
    .B2(_0661_),
    .X(_0452_));
 sky130_fd_sc_hd__mux2_1 _1164_ (.A0(\reg_temp[94] ),
    .A1(\reg_temp[12] ),
    .S(net585),
    .X(_0662_));
 sky130_fd_sc_hd__a22o_1 _1165_ (.A1(net1298),
    .A2(net529),
    .B1(net554),
    .B2(_0662_),
    .X(_0451_));
 sky130_fd_sc_hd__mux2_1 _1166_ (.A0(net1649),
    .A1(\reg_temp[11] ),
    .S(net585),
    .X(_0663_));
 sky130_fd_sc_hd__a22o_1 _1167_ (.A1(net1286),
    .A2(net529),
    .B1(net554),
    .B2(_0663_),
    .X(_0450_));
 sky130_fd_sc_hd__mux2_1 _1168_ (.A0(net1645),
    .A1(\reg_temp[10] ),
    .S(net585),
    .X(_0664_));
 sky130_fd_sc_hd__a22o_1 _1169_ (.A1(net1284),
    .A2(net529),
    .B1(net554),
    .B2(_0664_),
    .X(_0449_));
 sky130_fd_sc_hd__mux2_1 _1170_ (.A0(\reg_temp[91] ),
    .A1(\reg_temp[9] ),
    .S(net585),
    .X(_0665_));
 sky130_fd_sc_hd__a22o_1 _1171_ (.A1(net1281),
    .A2(net527),
    .B1(net552),
    .B2(_0665_),
    .X(_0448_));
 sky130_fd_sc_hd__mux2_1 _1172_ (.A0(\reg_temp[90] ),
    .A1(\reg_temp[8] ),
    .S(net585),
    .X(_0666_));
 sky130_fd_sc_hd__a22o_1 _1173_ (.A1(net1295),
    .A2(net529),
    .B1(net554),
    .B2(_0666_),
    .X(_0447_));
 sky130_fd_sc_hd__mux2_1 _1174_ (.A0(\reg_temp[89] ),
    .A1(\reg_temp[7] ),
    .S(net586),
    .X(_0667_));
 sky130_fd_sc_hd__a22o_1 _1175_ (.A1(net1280),
    .A2(net527),
    .B1(net552),
    .B2(_0667_),
    .X(_0446_));
 sky130_fd_sc_hd__mux2_1 _1176_ (.A0(\reg_temp[88] ),
    .A1(\reg_temp[6] ),
    .S(net586),
    .X(_0668_));
 sky130_fd_sc_hd__a22o_1 _1177_ (.A1(net1315),
    .A2(net529),
    .B1(net554),
    .B2(_0668_),
    .X(_0445_));
 sky130_fd_sc_hd__mux2_1 _1178_ (.A0(\reg_temp[87] ),
    .A1(\reg_temp[5] ),
    .S(net586),
    .X(_0669_));
 sky130_fd_sc_hd__a22o_1 _1179_ (.A1(net1261),
    .A2(net527),
    .B1(net552),
    .B2(_0669_),
    .X(_0444_));
 sky130_fd_sc_hd__mux2_1 _1180_ (.A0(net1636),
    .A1(net1640),
    .S(net585),
    .X(_0670_));
 sky130_fd_sc_hd__a22o_1 _1181_ (.A1(net1285),
    .A2(net529),
    .B1(net554),
    .B2(_0670_),
    .X(_0443_));
 sky130_fd_sc_hd__mux2_1 _1182_ (.A0(net1641),
    .A1(\reg_temp[3] ),
    .S(net585),
    .X(_0671_));
 sky130_fd_sc_hd__a22o_1 _1183_ (.A1(net1282),
    .A2(net529),
    .B1(net554),
    .B2(_0671_),
    .X(_0442_));
 sky130_fd_sc_hd__mux2_1 _1184_ (.A0(\reg_temp[84] ),
    .A1(\reg_temp[2] ),
    .S(net585),
    .X(_0672_));
 sky130_fd_sc_hd__a22o_1 _1185_ (.A1(net1260),
    .A2(net527),
    .B1(net552),
    .B2(_0672_),
    .X(_0441_));
 sky130_fd_sc_hd__mux2_1 _1186_ (.A0(\reg_temp[83] ),
    .A1(\reg_temp[1] ),
    .S(net585),
    .X(_0673_));
 sky130_fd_sc_hd__a22o_1 _1187_ (.A1(net1312),
    .A2(net527),
    .B1(net552),
    .B2(_0673_),
    .X(_0440_));
 sky130_fd_sc_hd__mux2_1 _1188_ (.A0(net1628),
    .A1(\reg_temp[0] ),
    .S(net585),
    .X(_0674_));
 sky130_fd_sc_hd__a22o_1 _1189_ (.A1(net1262),
    .A2(net527),
    .B1(net552),
    .B2(_0674_),
    .X(_0439_));
 sky130_fd_sc_hd__o21a_1 _1190_ (.A1(_0524_),
    .A2(net1151),
    .B1(net520),
    .X(_0675_));
 sky130_fd_sc_hd__or3_1 _1191_ (.A(net695),
    .B(net1219),
    .C(net1152),
    .X(_0438_));
 sky130_fd_sc_hd__and3b_1 _1192_ (.A_N(net1211),
    .B(_0564_),
    .C(net1200),
    .X(_0676_));
 sky130_fd_sc_hd__nand2_4 _1193_ (.A(_0524_),
    .B(_0570_),
    .Y(_0006_));
 sky130_fd_sc_hd__or3b_1 _1194_ (.A(_0576_),
    .B(net1212),
    .C_N(_0006_),
    .X(_0677_));
 sky130_fd_sc_hd__mux2_1 _1195_ (.A0(net695),
    .A1(net518),
    .S(net1213),
    .X(_0437_));
 sky130_fd_sc_hd__a21o_1 _1196_ (.A1(net517),
    .A2(net1213),
    .B1(net1206),
    .X(_0436_));
 sky130_fd_sc_hd__or4_1 _1197_ (.A(_0535_),
    .B(_0548_),
    .C(_0556_),
    .D(net564),
    .X(_0678_));
 sky130_fd_sc_hd__and3_1 _1198_ (.A(net560),
    .B(_0590_),
    .C(net778),
    .X(_0679_));
 sky130_fd_sc_hd__a21bo_1 _1199_ (.A1(net659),
    .A2(_0679_),
    .B1_N(_0678_),
    .X(_0680_));
 sky130_fd_sc_hd__mux2_1 _1200_ (.A0(net660),
    .A1(net516),
    .S(net1213),
    .X(_0435_));
 sky130_fd_sc_hd__and2_4 _1201_ (.A(\current_state[0] ),
    .B(\current_state[1] ),
    .X(_0007_));
 sky130_fd_sc_hd__a21oi_1 _1202_ (.A1(\current_state[0] ),
    .A2(net260),
    .B1(_0006_),
    .Y(_0681_));
 sky130_fd_sc_hd__a31o_1 _1203_ (.A1(_0552_),
    .A2(_0564_),
    .A3(net680),
    .B1(_0681_),
    .X(_0682_));
 sky130_fd_sc_hd__or3_1 _1204_ (.A(net695),
    .B(_0585_),
    .C(net681),
    .X(_0683_));
 sky130_fd_sc_hd__and2_1 _1205_ (.A(net595),
    .B(net927),
    .X(_0684_));
 sky130_fd_sc_hd__a21o_1 _1206_ (.A1(net70),
    .A2(net564),
    .B1(net928),
    .X(_0685_));
 sky130_fd_sc_hd__mux2_1 _1207_ (.A0(net929),
    .A1(\reg_temp[162] ),
    .S(net525),
    .X(_0434_));
 sky130_fd_sc_hd__and2_1 _1208_ (.A(net595),
    .B(net825),
    .X(_0686_));
 sky130_fd_sc_hd__a221o_1 _1209_ (.A1(net69),
    .A2(net570),
    .B1(net583),
    .B2(\reg_temp[162] ),
    .C1(net826),
    .X(_0687_));
 sky130_fd_sc_hd__mux2_1 _1210_ (.A0(_0687_),
    .A1(\reg_temp[161] ),
    .S(net525),
    .X(_0433_));
 sky130_fd_sc_hd__and2_1 _1211_ (.A(net595),
    .B(net887),
    .X(_0688_));
 sky130_fd_sc_hd__a221o_1 _1212_ (.A1(net68),
    .A2(net570),
    .B1(net583),
    .B2(\reg_temp[161] ),
    .C1(net888),
    .X(_0689_));
 sky130_fd_sc_hd__mux2_1 _1213_ (.A0(_0689_),
    .A1(\reg_temp[160] ),
    .S(net525),
    .X(_0432_));
 sky130_fd_sc_hd__and2_1 _1214_ (.A(net595),
    .B(net954),
    .X(_0690_));
 sky130_fd_sc_hd__a221o_1 _1215_ (.A1(net66),
    .A2(net569),
    .B1(net582),
    .B2(\reg_temp[160] ),
    .C1(net955),
    .X(_0691_));
 sky130_fd_sc_hd__mux2_1 _1216_ (.A0(_0691_),
    .A1(\reg_temp[159] ),
    .S(net525),
    .X(_0431_));
 sky130_fd_sc_hd__and2_1 _1217_ (.A(net595),
    .B(net1071),
    .X(_0692_));
 sky130_fd_sc_hd__a221o_1 _1218_ (.A1(net65),
    .A2(net568),
    .B1(net581),
    .B2(\reg_temp[159] ),
    .C1(net1072),
    .X(_0693_));
 sky130_fd_sc_hd__mux2_1 _1219_ (.A0(net1073),
    .A1(\reg_temp[158] ),
    .S(net525),
    .X(_0430_));
 sky130_fd_sc_hd__and2_1 _1220_ (.A(net595),
    .B(net1171),
    .X(_0694_));
 sky130_fd_sc_hd__a221o_1 _1221_ (.A1(net64),
    .A2(net568),
    .B1(net581),
    .B2(\reg_temp[158] ),
    .C1(net1172),
    .X(_0695_));
 sky130_fd_sc_hd__mux2_1 _1222_ (.A0(_0695_),
    .A1(\reg_temp[157] ),
    .S(net525),
    .X(_0429_));
 sky130_fd_sc_hd__and2_1 _1223_ (.A(net595),
    .B(net1099),
    .X(_0696_));
 sky130_fd_sc_hd__a221o_1 _1224_ (.A1(net63),
    .A2(net568),
    .B1(net581),
    .B2(\reg_temp[157] ),
    .C1(net1100),
    .X(_0697_));
 sky130_fd_sc_hd__mux2_1 _1225_ (.A0(net1101),
    .A1(\reg_temp[156] ),
    .S(net525),
    .X(_0428_));
 sky130_fd_sc_hd__and2_1 _1226_ (.A(net595),
    .B(net1078),
    .X(_0698_));
 sky130_fd_sc_hd__a221o_1 _1227_ (.A1(net62),
    .A2(net568),
    .B1(net581),
    .B2(\reg_temp[156] ),
    .C1(net1079),
    .X(_0699_));
 sky130_fd_sc_hd__mux2_1 _1228_ (.A0(_0699_),
    .A1(\reg_temp[155] ),
    .S(net525),
    .X(_0427_));
 sky130_fd_sc_hd__and2_1 _1229_ (.A(net595),
    .B(net1004),
    .X(_0700_));
 sky130_fd_sc_hd__a221o_1 _1230_ (.A1(net61),
    .A2(net568),
    .B1(net581),
    .B2(\reg_temp[155] ),
    .C1(net1005),
    .X(_0701_));
 sky130_fd_sc_hd__mux2_1 _1231_ (.A0(_0701_),
    .A1(\reg_temp[154] ),
    .S(net525),
    .X(_0426_));
 sky130_fd_sc_hd__and2_1 _1232_ (.A(net596),
    .B(net1040),
    .X(_0702_));
 sky130_fd_sc_hd__a221o_1 _1233_ (.A1(net60),
    .A2(net568),
    .B1(net581),
    .B2(\reg_temp[154] ),
    .C1(net1041),
    .X(_0703_));
 sky130_fd_sc_hd__mux2_1 _1234_ (.A0(_0703_),
    .A1(\reg_temp[153] ),
    .S(net525),
    .X(_0425_));
 sky130_fd_sc_hd__and2_1 _1235_ (.A(net596),
    .B(net1066),
    .X(_0704_));
 sky130_fd_sc_hd__a221o_1 _1236_ (.A1(net59),
    .A2(net569),
    .B1(net582),
    .B2(\reg_temp[153] ),
    .C1(net1067),
    .X(_0705_));
 sky130_fd_sc_hd__mux2_1 _1237_ (.A0(_0705_),
    .A1(\reg_temp[152] ),
    .S(net525),
    .X(_0424_));
 sky130_fd_sc_hd__and2_1 _1238_ (.A(net596),
    .B(net1092),
    .X(_0706_));
 sky130_fd_sc_hd__a221o_1 _1239_ (.A1(net58),
    .A2(net569),
    .B1(net582),
    .B2(\reg_temp[152] ),
    .C1(net1093),
    .X(_0707_));
 sky130_fd_sc_hd__mux2_1 _1240_ (.A0(_0707_),
    .A1(\reg_temp[151] ),
    .S(net525),
    .X(_0423_));
 sky130_fd_sc_hd__and2_1 _1241_ (.A(net596),
    .B(net1015),
    .X(_0708_));
 sky130_fd_sc_hd__a221o_1 _1242_ (.A1(net57),
    .A2(net569),
    .B1(net582),
    .B2(\reg_temp[151] ),
    .C1(net1016),
    .X(_0709_));
 sky130_fd_sc_hd__mux2_1 _1243_ (.A0(net1017),
    .A1(\reg_temp[150] ),
    .S(net525),
    .X(_0422_));
 sky130_fd_sc_hd__and2_1 _1244_ (.A(net596),
    .B(net1035),
    .X(_0710_));
 sky130_fd_sc_hd__a221o_1 _1245_ (.A1(net55),
    .A2(net570),
    .B1(net583),
    .B2(\reg_temp[150] ),
    .C1(net1036),
    .X(_0711_));
 sky130_fd_sc_hd__mux2_1 _1246_ (.A0(_0711_),
    .A1(\reg_temp[149] ),
    .S(net525),
    .X(_0421_));
 sky130_fd_sc_hd__and2_1 _1247_ (.A(net596),
    .B(net968),
    .X(_0712_));
 sky130_fd_sc_hd__a221o_1 _1248_ (.A1(net54),
    .A2(net570),
    .B1(net583),
    .B2(\reg_temp[149] ),
    .C1(net969),
    .X(_0713_));
 sky130_fd_sc_hd__mux2_1 _1249_ (.A0(net970),
    .A1(\reg_temp[148] ),
    .S(net525),
    .X(_0420_));
 sky130_fd_sc_hd__and2_1 _1250_ (.A(net596),
    .B(net981),
    .X(_0714_));
 sky130_fd_sc_hd__a221o_1 _1251_ (.A1(net53),
    .A2(net569),
    .B1(net582),
    .B2(\reg_temp[148] ),
    .C1(net982),
    .X(_0715_));
 sky130_fd_sc_hd__mux2_1 _1252_ (.A0(net983),
    .A1(\reg_temp[147] ),
    .S(net525),
    .X(_0419_));
 sky130_fd_sc_hd__and2_1 _1253_ (.A(net596),
    .B(net973),
    .X(_0716_));
 sky130_fd_sc_hd__a221o_1 _1254_ (.A1(net52),
    .A2(net568),
    .B1(net581),
    .B2(\reg_temp[147] ),
    .C1(net974),
    .X(_0717_));
 sky130_fd_sc_hd__mux2_1 _1255_ (.A0(net975),
    .A1(net1561),
    .S(net683),
    .X(_0418_));
 sky130_fd_sc_hd__and2_1 _1256_ (.A(net595),
    .B(net1131),
    .X(_0718_));
 sky130_fd_sc_hd__a221o_1 _1257_ (.A1(net51),
    .A2(net571),
    .B1(net584),
    .B2(\reg_temp[146] ),
    .C1(net1132),
    .X(_0719_));
 sky130_fd_sc_hd__mux2_1 _1258_ (.A0(_0719_),
    .A1(\reg_temp[145] ),
    .S(net683),
    .X(_0417_));
 sky130_fd_sc_hd__and2_1 _1259_ (.A(net595),
    .B(net963),
    .X(_0720_));
 sky130_fd_sc_hd__a221o_1 _1260_ (.A1(net50),
    .A2(net571),
    .B1(net584),
    .B2(\reg_temp[145] ),
    .C1(net964),
    .X(_0721_));
 sky130_fd_sc_hd__mux2_1 _1261_ (.A0(_0721_),
    .A1(\reg_temp[144] ),
    .S(net683),
    .X(_0416_));
 sky130_fd_sc_hd__and2_1 _1262_ (.A(net595),
    .B(net1029),
    .X(_0722_));
 sky130_fd_sc_hd__a221o_1 _1263_ (.A1(net49),
    .A2(net571),
    .B1(net584),
    .B2(\reg_temp[144] ),
    .C1(net1030),
    .X(_0723_));
 sky130_fd_sc_hd__mux2_1 _1264_ (.A0(net1031),
    .A1(net1581),
    .S(net683),
    .X(_0415_));
 sky130_fd_sc_hd__and2_1 _1265_ (.A(net596),
    .B(net1156),
    .X(_0724_));
 sky130_fd_sc_hd__a221o_1 _1266_ (.A1(net48),
    .A2(net571),
    .B1(net584),
    .B2(\reg_temp[143] ),
    .C1(net1157),
    .X(_0725_));
 sky130_fd_sc_hd__mux2_1 _1267_ (.A0(net1158),
    .A1(\reg_temp[142] ),
    .S(net683),
    .X(_0414_));
 sky130_fd_sc_hd__and2_1 _1268_ (.A(net596),
    .B(net1119),
    .X(_0726_));
 sky130_fd_sc_hd__a221o_1 _1269_ (.A1(net47),
    .A2(net571),
    .B1(net584),
    .B2(\reg_temp[142] ),
    .C1(net1120),
    .X(_0727_));
 sky130_fd_sc_hd__mux2_1 _1270_ (.A0(_0727_),
    .A1(\reg_temp[141] ),
    .S(net524),
    .X(_0413_));
 sky130_fd_sc_hd__and2_1 _1271_ (.A(net596),
    .B(net1126),
    .X(_0728_));
 sky130_fd_sc_hd__a221o_1 _1272_ (.A1(net46),
    .A2(net571),
    .B1(net584),
    .B2(\reg_temp[141] ),
    .C1(net1127),
    .X(_0729_));
 sky130_fd_sc_hd__mux2_1 _1273_ (.A0(_0729_),
    .A1(\reg_temp[140] ),
    .S(net524),
    .X(_0412_));
 sky130_fd_sc_hd__and2_1 _1274_ (.A(net595),
    .B(net996),
    .X(_0730_));
 sky130_fd_sc_hd__a221o_1 _1275_ (.A1(net44),
    .A2(net566),
    .B1(net579),
    .B2(\reg_temp[140] ),
    .C1(net997),
    .X(_0731_));
 sky130_fd_sc_hd__mux2_1 _1276_ (.A0(net998),
    .A1(net1631),
    .S(net524),
    .X(_0411_));
 sky130_fd_sc_hd__and2_1 _1277_ (.A(net595),
    .B(net1106),
    .X(_0732_));
 sky130_fd_sc_hd__a221o_1 _1278_ (.A1(net43),
    .A2(net571),
    .B1(net584),
    .B2(\reg_temp[139] ),
    .C1(net1107),
    .X(_0733_));
 sky130_fd_sc_hd__mux2_1 _1279_ (.A0(net1108),
    .A1(net1614),
    .S(net524),
    .X(_0410_));
 sky130_fd_sc_hd__and2_1 _1280_ (.A(net597),
    .B(net1047),
    .X(_0734_));
 sky130_fd_sc_hd__a221o_1 _1281_ (.A1(net42),
    .A2(net567),
    .B1(net580),
    .B2(\reg_temp[138] ),
    .C1(net1048),
    .X(_0735_));
 sky130_fd_sc_hd__mux2_1 _1282_ (.A0(_0735_),
    .A1(\reg_temp[137] ),
    .S(net683),
    .X(_0409_));
 sky130_fd_sc_hd__and2_1 _1283_ (.A(net597),
    .B(net1057),
    .X(_0736_));
 sky130_fd_sc_hd__a221o_1 _1284_ (.A1(net41),
    .A2(net566),
    .B1(net579),
    .B2(\reg_temp[137] ),
    .C1(net1058),
    .X(_0737_));
 sky130_fd_sc_hd__mux2_1 _1285_ (.A0(_0737_),
    .A1(\reg_temp[136] ),
    .S(net524),
    .X(_0408_));
 sky130_fd_sc_hd__and2_1 _1286_ (.A(net597),
    .B(net1009),
    .X(_0738_));
 sky130_fd_sc_hd__a221o_1 _1287_ (.A1(net40),
    .A2(net566),
    .B1(net579),
    .B2(\reg_temp[136] ),
    .C1(net1010),
    .X(_0739_));
 sky130_fd_sc_hd__mux2_1 _1288_ (.A0(net1011),
    .A1(\reg_temp[135] ),
    .S(net524),
    .X(_0407_));
 sky130_fd_sc_hd__and2_1 _1289_ (.A(net597),
    .B(net941),
    .X(_0740_));
 sky130_fd_sc_hd__a221o_1 _1290_ (.A1(net39),
    .A2(net566),
    .B1(net579),
    .B2(\reg_temp[135] ),
    .C1(net942),
    .X(_0741_));
 sky130_fd_sc_hd__mux2_1 _1291_ (.A0(net943),
    .A1(\reg_temp[134] ),
    .S(net524),
    .X(_0406_));
 sky130_fd_sc_hd__and2_1 _1292_ (.A(net597),
    .B(net922),
    .X(_0742_));
 sky130_fd_sc_hd__a221o_1 _1293_ (.A1(net38),
    .A2(net566),
    .B1(net579),
    .B2(\reg_temp[134] ),
    .C1(net923),
    .X(_0743_));
 sky130_fd_sc_hd__mux2_1 _1294_ (.A0(net924),
    .A1(\reg_temp[133] ),
    .S(net524),
    .X(_0405_));
 sky130_fd_sc_hd__and2_1 _1295_ (.A(net597),
    .B(net820),
    .X(_0744_));
 sky130_fd_sc_hd__a221o_1 _1296_ (.A1(net37),
    .A2(net566),
    .B1(net579),
    .B2(\reg_temp[133] ),
    .C1(net821),
    .X(_0745_));
 sky130_fd_sc_hd__mux2_1 _1297_ (.A0(net822),
    .A1(\reg_temp[132] ),
    .S(net524),
    .X(_0404_));
 sky130_fd_sc_hd__and2_1 _1298_ (.A(net597),
    .B(net803),
    .X(_0746_));
 sky130_fd_sc_hd__a221o_1 _1299_ (.A1(net36),
    .A2(net566),
    .B1(net579),
    .B2(\reg_temp[132] ),
    .C1(net804),
    .X(_0747_));
 sky130_fd_sc_hd__mux2_1 _1300_ (.A0(_0747_),
    .A1(\reg_temp[131] ),
    .S(net524),
    .X(_0403_));
 sky130_fd_sc_hd__and2_1 _1301_ (.A(net597),
    .B(net797),
    .X(_0748_));
 sky130_fd_sc_hd__a221o_1 _1302_ (.A1(net35),
    .A2(net564),
    .B1(net580),
    .B2(\reg_temp[131] ),
    .C1(net798),
    .X(_0749_));
 sky130_fd_sc_hd__mux2_1 _1303_ (.A0(net799),
    .A1(\reg_temp[130] ),
    .S(net524),
    .X(_0402_));
 sky130_fd_sc_hd__and2_1 _1304_ (.A(net597),
    .B(net751),
    .X(_0750_));
 sky130_fd_sc_hd__a221o_1 _1305_ (.A1(net33),
    .A2(net567),
    .B1(net577),
    .B2(\reg_temp[130] ),
    .C1(net752),
    .X(_0751_));
 sky130_fd_sc_hd__mux2_1 _1306_ (.A0(net753),
    .A1(\reg_temp[129] ),
    .S(net524),
    .X(_0401_));
 sky130_fd_sc_hd__and2_1 _1307_ (.A(net597),
    .B(net715),
    .X(_0752_));
 sky130_fd_sc_hd__a221o_1 _1308_ (.A1(net32),
    .A2(net564),
    .B1(net577),
    .B2(\reg_temp[129] ),
    .C1(net716),
    .X(_0753_));
 sky130_fd_sc_hd__mux2_1 _1309_ (.A0(net717),
    .A1(\reg_temp[128] ),
    .S(net524),
    .X(_0400_));
 sky130_fd_sc_hd__and2_1 _1310_ (.A(net597),
    .B(net668),
    .X(_0754_));
 sky130_fd_sc_hd__a221o_1 _1311_ (.A1(net31),
    .A2(net564),
    .B1(net577),
    .B2(\reg_temp[128] ),
    .C1(net669),
    .X(_0755_));
 sky130_fd_sc_hd__mux2_1 _1312_ (.A0(net670),
    .A1(\reg_temp[127] ),
    .S(net524),
    .X(_0399_));
 sky130_fd_sc_hd__and2_1 _1313_ (.A(net593),
    .B(net853),
    .X(_0756_));
 sky130_fd_sc_hd__a221o_1 _1314_ (.A1(net30),
    .A2(net564),
    .B1(net580),
    .B2(\reg_temp[127] ),
    .C1(net854),
    .X(_0757_));
 sky130_fd_sc_hd__mux2_1 _1315_ (.A0(net855),
    .A1(net1588),
    .S(net524),
    .X(_0398_));
 sky130_fd_sc_hd__and2_1 _1316_ (.A(net593),
    .B(net700),
    .X(_0758_));
 sky130_fd_sc_hd__a221o_1 _1317_ (.A1(net29),
    .A2(net567),
    .B1(net577),
    .B2(\reg_temp[126] ),
    .C1(net701),
    .X(_0759_));
 sky130_fd_sc_hd__mux2_1 _1318_ (.A0(net702),
    .A1(\reg_temp[125] ),
    .S(net524),
    .X(_0397_));
 sky130_fd_sc_hd__and2_1 _1319_ (.A(net593),
    .B(net728),
    .X(_0760_));
 sky130_fd_sc_hd__a221o_1 _1320_ (.A1(net28),
    .A2(net567),
    .B1(net577),
    .B2(\reg_temp[125] ),
    .C1(net729),
    .X(_0761_));
 sky130_fd_sc_hd__mux2_1 _1321_ (.A0(net730),
    .A1(\reg_temp[124] ),
    .S(net684),
    .X(_0396_));
 sky130_fd_sc_hd__and2_1 _1322_ (.A(net593),
    .B(net839),
    .X(_0762_));
 sky130_fd_sc_hd__a221o_1 _1323_ (.A1(net27),
    .A2(net564),
    .B1(net577),
    .B2(\reg_temp[124] ),
    .C1(net840),
    .X(_0763_));
 sky130_fd_sc_hd__mux2_1 _1324_ (.A0(_0763_),
    .A1(\reg_temp[123] ),
    .S(net684),
    .X(_0395_));
 sky130_fd_sc_hd__and2_1 _1325_ (.A(net593),
    .B(net847),
    .X(_0764_));
 sky130_fd_sc_hd__a221o_1 _1326_ (.A1(net26),
    .A2(net564),
    .B1(net577),
    .B2(\reg_temp[123] ),
    .C1(net848),
    .X(_0765_));
 sky130_fd_sc_hd__mux2_1 _1327_ (.A0(_0765_),
    .A1(\reg_temp[122] ),
    .S(net684),
    .X(_0394_));
 sky130_fd_sc_hd__and2_1 _1328_ (.A(net593),
    .B(net910),
    .X(_0766_));
 sky130_fd_sc_hd__a221o_1 _1329_ (.A1(net25),
    .A2(net564),
    .B1(net577),
    .B2(\reg_temp[122] ),
    .C1(net911),
    .X(_0767_));
 sky130_fd_sc_hd__mux2_1 _1330_ (.A0(net912),
    .A1(net1618),
    .S(net684),
    .X(_0393_));
 sky130_fd_sc_hd__and2_1 _1331_ (.A(net593),
    .B(net883),
    .X(_0768_));
 sky130_fd_sc_hd__a221o_1 _1332_ (.A1(net24),
    .A2(net564),
    .B1(net577),
    .B2(\reg_temp[121] ),
    .C1(net884),
    .X(_0769_));
 sky130_fd_sc_hd__mux2_1 _1333_ (.A0(net885),
    .A1(net1605),
    .S(net684),
    .X(_0392_));
 sky130_fd_sc_hd__and2_1 _1334_ (.A(net593),
    .B(net992),
    .X(_0770_));
 sky130_fd_sc_hd__a221o_1 _1335_ (.A1(net22),
    .A2(net565),
    .B1(net578),
    .B2(\reg_temp[120] ),
    .C1(net993),
    .X(_0771_));
 sky130_fd_sc_hd__mux2_1 _1336_ (.A0(net994),
    .A1(net1625),
    .S(net684),
    .X(_0391_));
 sky130_fd_sc_hd__and2_1 _1337_ (.A(net593),
    .B(net1000),
    .X(_0772_));
 sky130_fd_sc_hd__a221o_1 _1338_ (.A1(net21),
    .A2(net565),
    .B1(net578),
    .B2(\reg_temp[119] ),
    .C1(net1001),
    .X(_0773_));
 sky130_fd_sc_hd__mux2_1 _1339_ (.A0(_0773_),
    .A1(\reg_temp[118] ),
    .S(net523),
    .X(_0390_));
 sky130_fd_sc_hd__and2_1 _1340_ (.A(net593),
    .B(net1025),
    .X(_0774_));
 sky130_fd_sc_hd__a221o_1 _1341_ (.A1(net20),
    .A2(net565),
    .B1(net578),
    .B2(\reg_temp[118] ),
    .C1(net1026),
    .X(_0775_));
 sky130_fd_sc_hd__mux2_1 _1342_ (.A0(_0775_),
    .A1(\reg_temp[117] ),
    .S(net523),
    .X(_0389_));
 sky130_fd_sc_hd__and2_1 _1343_ (.A(net592),
    .B(net792),
    .X(_0776_));
 sky130_fd_sc_hd__a221o_1 _1344_ (.A1(net19),
    .A2(net565),
    .B1(net578),
    .B2(\reg_temp[117] ),
    .C1(net793),
    .X(_0777_));
 sky130_fd_sc_hd__mux2_1 _1345_ (.A0(_0777_),
    .A1(net1592),
    .S(net522),
    .X(_0388_));
 sky130_fd_sc_hd__and2_1 _1346_ (.A(net592),
    .B(net762),
    .X(_0778_));
 sky130_fd_sc_hd__a221o_1 _1347_ (.A1(net18),
    .A2(net565),
    .B1(net578),
    .B2(\reg_temp[116] ),
    .C1(net763),
    .X(_0779_));
 sky130_fd_sc_hd__mux2_1 _1348_ (.A0(net764),
    .A1(net1635),
    .S(net523),
    .X(_0387_));
 sky130_fd_sc_hd__and2_1 _1349_ (.A(net593),
    .B(net1062),
    .X(_0780_));
 sky130_fd_sc_hd__a221o_1 _1350_ (.A1(net17),
    .A2(net565),
    .B1(net578),
    .B2(\reg_temp[115] ),
    .C1(net1063),
    .X(_0781_));
 sky130_fd_sc_hd__mux2_1 _1351_ (.A0(_0781_),
    .A1(net1616),
    .S(net522),
    .X(_0386_));
 sky130_fd_sc_hd__and2_1 _1352_ (.A(net592),
    .B(net900),
    .X(_0782_));
 sky130_fd_sc_hd__a221o_1 _1353_ (.A1(net16),
    .A2(net565),
    .B1(net579),
    .B2(\reg_temp[114] ),
    .C1(net901),
    .X(_0783_));
 sky130_fd_sc_hd__mux2_1 _1354_ (.A0(_0783_),
    .A1(net1598),
    .S(net523),
    .X(_0385_));
 sky130_fd_sc_hd__and2_1 _1355_ (.A(net592),
    .B(net932),
    .X(_0784_));
 sky130_fd_sc_hd__a221o_1 _1356_ (.A1(net15),
    .A2(net565),
    .B1(net579),
    .B2(\reg_temp[113] ),
    .C1(net933),
    .X(_0785_));
 sky130_fd_sc_hd__mux2_1 _1357_ (.A0(net934),
    .A1(net1601),
    .S(net523),
    .X(_0384_));
 sky130_fd_sc_hd__and2_1 _1358_ (.A(net592),
    .B(net946),
    .X(_0786_));
 sky130_fd_sc_hd__a221o_1 _1359_ (.A1(net14),
    .A2(net566),
    .B1(net579),
    .B2(\reg_temp[112] ),
    .C1(net947),
    .X(_0787_));
 sky130_fd_sc_hd__mux2_1 _1360_ (.A0(_0787_),
    .A1(\reg_temp[111] ),
    .S(net523),
    .X(_0383_));
 sky130_fd_sc_hd__and2_1 _1361_ (.A(net592),
    .B(net879),
    .X(_0788_));
 sky130_fd_sc_hd__a221o_1 _1362_ (.A1(net13),
    .A2(net566),
    .B1(net578),
    .B2(\reg_temp[111] ),
    .C1(net880),
    .X(_0789_));
 sky130_fd_sc_hd__mux2_1 _1363_ (.A0(_0789_),
    .A1(net1604),
    .S(net523),
    .X(_0382_));
 sky130_fd_sc_hd__and2_1 _1364_ (.A(net592),
    .B(net893),
    .X(_0790_));
 sky130_fd_sc_hd__a221o_1 _1365_ (.A1(net11),
    .A2(net566),
    .B1(net578),
    .B2(\reg_temp[110] ),
    .C1(net894),
    .X(_0791_));
 sky130_fd_sc_hd__mux2_1 _1366_ (.A0(_0791_),
    .A1(net1583),
    .S(net523),
    .X(_0381_));
 sky130_fd_sc_hd__and2_1 _1367_ (.A(net592),
    .B(net904),
    .X(_0792_));
 sky130_fd_sc_hd__a221o_1 _1368_ (.A1(net10),
    .A2(net566),
    .B1(net578),
    .B2(\reg_temp[109] ),
    .C1(net905),
    .X(_0793_));
 sky130_fd_sc_hd__mux2_1 _1369_ (.A0(net906),
    .A1(\reg_temp[108] ),
    .S(net523),
    .X(_0380_));
 sky130_fd_sc_hd__and2_1 _1370_ (.A(net592),
    .B(net864),
    .X(_0794_));
 sky130_fd_sc_hd__a221o_1 _1371_ (.A1(net9),
    .A2(net565),
    .B1(net578),
    .B2(\reg_temp[108] ),
    .C1(net865),
    .X(_0795_));
 sky130_fd_sc_hd__mux2_1 _1372_ (.A0(_0795_),
    .A1(\reg_temp[107] ),
    .S(net523),
    .X(_0379_));
 sky130_fd_sc_hd__and2_1 _1373_ (.A(net592),
    .B(net783),
    .X(_0796_));
 sky130_fd_sc_hd__a221o_1 _1374_ (.A1(net8),
    .A2(net565),
    .B1(net578),
    .B2(\reg_temp[107] ),
    .C1(net784),
    .X(_0797_));
 sky130_fd_sc_hd__mux2_1 _1375_ (.A0(net785),
    .A1(\reg_temp[106] ),
    .S(net522),
    .X(_0378_));
 sky130_fd_sc_hd__and2_1 _1376_ (.A(net594),
    .B(net1192),
    .X(_0798_));
 sky130_fd_sc_hd__a221o_1 _1377_ (.A1(net7),
    .A2(net565),
    .B1(net578),
    .B2(\reg_temp[106] ),
    .C1(net1193),
    .X(_0799_));
 sky130_fd_sc_hd__mux2_1 _1378_ (.A0(net1194),
    .A1(net1643),
    .S(net683),
    .X(_0377_));
 sky130_fd_sc_hd__and2_1 _1379_ (.A(net594),
    .B(net1181),
    .X(_0800_));
 sky130_fd_sc_hd__a221o_1 _1380_ (.A1(net6),
    .A2(net566),
    .B1(net579),
    .B2(\reg_temp[105] ),
    .C1(net1182),
    .X(_0801_));
 sky130_fd_sc_hd__mux2_1 _1381_ (.A0(_0801_),
    .A1(net1582),
    .S(net522),
    .X(_0376_));
 sky130_fd_sc_hd__and2_1 _1382_ (.A(net594),
    .B(net1185),
    .X(_0802_));
 sky130_fd_sc_hd__a221o_1 _1383_ (.A1(net5),
    .A2(net565),
    .B1(net578),
    .B2(\reg_temp[104] ),
    .C1(net1186),
    .X(_0803_));
 sky130_fd_sc_hd__mux2_1 _1384_ (.A0(_0803_),
    .A1(net1612),
    .S(net522),
    .X(_0375_));
 sky130_fd_sc_hd__and2_1 _1385_ (.A(net594),
    .B(net1177),
    .X(_0804_));
 sky130_fd_sc_hd__a221o_1 _1386_ (.A1(net4),
    .A2(net565),
    .B1(net579),
    .B2(\reg_temp[103] ),
    .C1(net1178),
    .X(_0805_));
 sky130_fd_sc_hd__mux2_1 _1387_ (.A0(net1179),
    .A1(net1632),
    .S(net522),
    .X(_0374_));
 sky130_fd_sc_hd__and2_2 _1388_ (.A(net594),
    .B(net659),
    .X(_0806_));
 sky130_fd_sc_hd__a221o_1 _1389_ (.A1(net3),
    .A2(net563),
    .B1(net576),
    .B2(\reg_temp[102] ),
    .C1(_0806_),
    .X(_0807_));
 sky130_fd_sc_hd__mux2_1 _1390_ (.A0(_0807_),
    .A1(net1623),
    .S(net522),
    .X(_0373_));
 sky130_fd_sc_hd__and2_2 _1391_ (.A(net594),
    .B(net745),
    .X(_0808_));
 sky130_fd_sc_hd__a221o_1 _1392_ (.A1(net2),
    .A2(net563),
    .B1(net576),
    .B2(\reg_temp[101] ),
    .C1(_0808_),
    .X(_0809_));
 sky130_fd_sc_hd__mux2_1 _1393_ (.A0(_0809_),
    .A1(net1627),
    .S(net522),
    .X(_0372_));
 sky130_fd_sc_hd__and2_1 _1394_ (.A(net594),
    .B(net777),
    .X(_0810_));
 sky130_fd_sc_hd__a221o_1 _1395_ (.A1(net162),
    .A2(net563),
    .B1(net576),
    .B2(\reg_temp[100] ),
    .C1(_0810_),
    .X(_0811_));
 sky130_fd_sc_hd__mux2_1 _1396_ (.A0(_0811_),
    .A1(net1579),
    .S(net522),
    .X(_0371_));
 sky130_fd_sc_hd__nor2_1 _1397_ (.A(\current_state[1] ),
    .B(net1168),
    .Y(_0812_));
 sky130_fd_sc_hd__a221o_1 _1398_ (.A1(net161),
    .A2(net566),
    .B1(net579),
    .B2(\reg_temp[99] ),
    .C1(net1169),
    .X(_0813_));
 sky130_fd_sc_hd__mux2_1 _1399_ (.A0(_0813_),
    .A1(net1432),
    .S(net522),
    .X(_0370_));
 sky130_fd_sc_hd__and2_1 _1400_ (.A(net592),
    .B(net788),
    .X(_0814_));
 sky130_fd_sc_hd__a221o_1 _1401_ (.A1(net160),
    .A2(net565),
    .B1(net578),
    .B2(\reg_temp[98] ),
    .C1(net789),
    .X(_0815_));
 sky130_fd_sc_hd__mux2_1 _1402_ (.A0(net790),
    .A1(net1580),
    .S(net522),
    .X(_0369_));
 sky130_fd_sc_hd__and2_1 _1403_ (.A(net592),
    .B(net741),
    .X(_0816_));
 sky130_fd_sc_hd__a221o_1 _1404_ (.A1(net159),
    .A2(net563),
    .B1(net576),
    .B2(\reg_temp[97] ),
    .C1(net742),
    .X(_0817_));
 sky130_fd_sc_hd__mux2_1 _1405_ (.A0(net743),
    .A1(net1606),
    .S(net522),
    .X(_0368_));
 sky130_fd_sc_hd__and2_1 _1406_ (.A(net592),
    .B(net875),
    .X(_0818_));
 sky130_fd_sc_hd__a221o_1 _1407_ (.A1(net158),
    .A2(_0569_),
    .B1(net576),
    .B2(\reg_temp[96] ),
    .C1(net876),
    .X(_0819_));
 sky130_fd_sc_hd__mux2_1 _1408_ (.A0(_0819_),
    .A1(net1610),
    .S(net684),
    .X(_0367_));
 sky130_fd_sc_hd__and2_1 _1409_ (.A(net592),
    .B(net859),
    .X(_0820_));
 sky130_fd_sc_hd__a221o_1 _1410_ (.A1(net157),
    .A2(net563),
    .B1(_0007_),
    .B2(\reg_temp[95] ),
    .C1(net860),
    .X(_0821_));
 sky130_fd_sc_hd__mux2_1 _1411_ (.A0(_0821_),
    .A1(\reg_temp[94] ),
    .S(net684),
    .X(_0366_));
 sky130_fd_sc_hd__and2_1 _1412_ (.A(net592),
    .B(net812),
    .X(_0822_));
 sky130_fd_sc_hd__a221o_1 _1413_ (.A1(net156),
    .A2(net560),
    .B1(net573),
    .B2(\reg_temp[94] ),
    .C1(net813),
    .X(_0823_));
 sky130_fd_sc_hd__mux2_1 _1414_ (.A0(_0823_),
    .A1(\reg_temp[93] ),
    .S(net684),
    .X(_0365_));
 sky130_fd_sc_hd__and2_1 _1415_ (.A(net592),
    .B(net710),
    .X(_0824_));
 sky130_fd_sc_hd__a221o_1 _1416_ (.A1(net155),
    .A2(net559),
    .B1(net573),
    .B2(\reg_temp[93] ),
    .C1(net711),
    .X(_0825_));
 sky130_fd_sc_hd__mux2_1 _1417_ (.A0(_0825_),
    .A1(\reg_temp[92] ),
    .S(net684),
    .X(_0364_));
 sky130_fd_sc_hd__and2_1 _1418_ (.A(net591),
    .B(net757),
    .X(_0826_));
 sky130_fd_sc_hd__a221o_1 _1419_ (.A1(net154),
    .A2(net560),
    .B1(net573),
    .B2(\reg_temp[92] ),
    .C1(net758),
    .X(_0827_));
 sky130_fd_sc_hd__mux2_1 _1420_ (.A0(_0827_),
    .A1(\reg_temp[91] ),
    .S(net684),
    .X(_0363_));
 sky130_fd_sc_hd__and2_1 _1421_ (.A(net591),
    .B(net843),
    .X(_0828_));
 sky130_fd_sc_hd__a221o_1 _1422_ (.A1(net153),
    .A2(net563),
    .B1(net576),
    .B2(\reg_temp[91] ),
    .C1(net844),
    .X(_0829_));
 sky130_fd_sc_hd__mux2_1 _1423_ (.A0(_0829_),
    .A1(\reg_temp[90] ),
    .S(net684),
    .X(_0362_));
 sky130_fd_sc_hd__and2_1 _1424_ (.A(net591),
    .B(net773),
    .X(_0830_));
 sky130_fd_sc_hd__a221o_1 _1425_ (.A1(net151),
    .A2(net563),
    .B1(net576),
    .B2(\reg_temp[90] ),
    .C1(net774),
    .X(_0831_));
 sky130_fd_sc_hd__mux2_1 _1426_ (.A0(net775),
    .A1(net1634),
    .S(net522),
    .X(_0361_));
 sky130_fd_sc_hd__and2_1 _1427_ (.A(net591),
    .B(net720),
    .X(_0832_));
 sky130_fd_sc_hd__a221o_1 _1428_ (.A1(net150),
    .A2(net563),
    .B1(net576),
    .B2(\reg_temp[89] ),
    .C1(net721),
    .X(_0833_));
 sky130_fd_sc_hd__mux2_1 _1429_ (.A0(net722),
    .A1(\reg_temp[88] ),
    .S(net522),
    .X(_0360_));
 sky130_fd_sc_hd__and2_1 _1430_ (.A(net591),
    .B(net724),
    .X(_0834_));
 sky130_fd_sc_hd__a221o_1 _1431_ (.A1(net149),
    .A2(net563),
    .B1(net576),
    .B2(\reg_temp[88] ),
    .C1(net725),
    .X(_0835_));
 sky130_fd_sc_hd__mux2_1 _1432_ (.A0(net726),
    .A1(net1624),
    .S(net522),
    .X(_0359_));
 sky130_fd_sc_hd__and2_1 _1433_ (.A(net591),
    .B(net937),
    .X(_0836_));
 sky130_fd_sc_hd__a221o_1 _1434_ (.A1(net148),
    .A2(net563),
    .B1(net576),
    .B2(\reg_temp[87] ),
    .C1(net938),
    .X(_0837_));
 sky130_fd_sc_hd__mux2_1 _1435_ (.A0(net939),
    .A1(net1636),
    .S(net522),
    .X(_0358_));
 sky130_fd_sc_hd__and2_1 _1436_ (.A(net591),
    .B(net832),
    .X(_0838_));
 sky130_fd_sc_hd__a221o_1 _1437_ (.A1(net147),
    .A2(net560),
    .B1(net573),
    .B2(\reg_temp[86] ),
    .C1(net833),
    .X(_0839_));
 sky130_fd_sc_hd__mux2_1 _1438_ (.A0(_0839_),
    .A1(\reg_temp[85] ),
    .S(net684),
    .X(_0357_));
 sky130_fd_sc_hd__and2_1 _1439_ (.A(net591),
    .B(net673),
    .X(_0840_));
 sky130_fd_sc_hd__a221o_1 _1440_ (.A1(net146),
    .A2(net559),
    .B1(net573),
    .B2(\reg_temp[85] ),
    .C1(net674),
    .X(_0841_));
 sky130_fd_sc_hd__mux2_1 _1441_ (.A0(_0841_),
    .A1(\reg_temp[84] ),
    .S(net684),
    .X(_0356_));
 sky130_fd_sc_hd__and2_1 _1442_ (.A(net591),
    .B(net687),
    .X(_0842_));
 sky130_fd_sc_hd__a221o_1 _1443_ (.A1(net145),
    .A2(net560),
    .B1(net573),
    .B2(\reg_temp[84] ),
    .C1(net688),
    .X(_0843_));
 sky130_fd_sc_hd__mux2_1 _1444_ (.A0(_0843_),
    .A1(\reg_temp[83] ),
    .S(net684),
    .X(_0355_));
 sky130_fd_sc_hd__and2_1 _1445_ (.A(net591),
    .B(net705),
    .X(_0844_));
 sky130_fd_sc_hd__a221o_1 _1446_ (.A1(net144),
    .A2(net560),
    .B1(net573),
    .B2(\reg_temp[83] ),
    .C1(net706),
    .X(_0845_));
 sky130_fd_sc_hd__mux2_1 _1447_ (.A0(_0845_),
    .A1(\reg_temp[82] ),
    .S(net684),
    .X(_0354_));
 sky130_fd_sc_hd__a21bo_2 _1448_ (.A1(net1200),
    .A2(net735),
    .B1_N(_0574_),
    .X(_0846_));
 sky130_fd_sc_hd__mux2_1 _1449_ (.A0(net1200),
    .A1(net444),
    .S(_0846_),
    .X(_0353_));
 sky130_fd_sc_hd__a31o_1 _1450_ (.A1(net659),
    .A2(net745),
    .A3(_0679_),
    .B1(net573),
    .X(_0847_));
 sky130_fd_sc_hd__a21o_1 _1451_ (.A1(_0540_),
    .A2(_0564_),
    .B1(net746),
    .X(_0848_));
 sky130_fd_sc_hd__mux2_1 _1452_ (.A0(net747),
    .A1(net443),
    .S(_0846_),
    .X(_0352_));
 sky130_fd_sc_hd__or4_1 _1453_ (.A(net1142),
    .B(net1084),
    .C(net250),
    .D(_0544_),
    .X(_0849_));
 sky130_fd_sc_hd__a31oi_1 _1454_ (.A1(_0520_),
    .A2(_0526_),
    .A3(_0554_),
    .B1(net679),
    .Y(_0850_));
 sky130_fd_sc_hd__and4_1 _1455_ (.A(_0523_),
    .B(_0532_),
    .C(net1143),
    .D(_0850_),
    .X(_0851_));
 sky130_fd_sc_hd__xor2_1 _1456_ (.A(net659),
    .B(net745),
    .X(_0852_));
 sky130_fd_sc_hd__a211o_1 _1457_ (.A1(_0679_),
    .A2(_0852_),
    .B1(net1144),
    .C1(net573),
    .X(_0853_));
 sky130_fd_sc_hd__mux2_1 _1458_ (.A0(net1145),
    .A1(net442),
    .S(_0846_),
    .X(_0351_));
 sky130_fd_sc_hd__a41oi_1 _1459_ (.A1(_0532_),
    .A2(_0537_),
    .A3(_0567_),
    .A4(net767),
    .B1(_0524_),
    .Y(_0854_));
 sky130_fd_sc_hd__a211o_1 _1460_ (.A1(net567),
    .A2(net779),
    .B1(net577),
    .C1(net768),
    .X(_0855_));
 sky130_fd_sc_hd__mux2_1 _1461_ (.A0(net780),
    .A1(net441),
    .S(_0846_),
    .X(_0350_));
 sky130_fd_sc_hd__a211o_1 _1462_ (.A1(net567),
    .A2(net779),
    .B1(net1088),
    .C1(net595),
    .X(_0856_));
 sky130_fd_sc_hd__and2_1 _1463_ (.A(\reg_temp[81] ),
    .B(net570),
    .X(_0857_));
 sky130_fd_sc_hd__mux2_1 _1464_ (.A0(_0857_),
    .A1(net440),
    .S(net1089),
    .X(_0349_));
 sky130_fd_sc_hd__a21bo_1 _1465_ (.A1(net1234),
    .A2(net1221),
    .B1_N(net532),
    .X(_0348_));
 sky130_fd_sc_hd__mux2_1 _1466_ (.A0(_0006_),
    .A1(net445),
    .S(net1221),
    .X(_0347_));
 sky130_fd_sc_hd__a211o_1 _1467_ (.A1(_0552_),
    .A2(net735),
    .B1(_0681_),
    .C1(net768),
    .X(_0858_));
 sky130_fd_sc_hd__a22o_1 _1468_ (.A1(net597),
    .A2(net663),
    .B1(net577),
    .B2(\reg_temp[82] ),
    .X(_0859_));
 sky130_fd_sc_hd__a21o_1 _1469_ (.A1(net143),
    .A2(net564),
    .B1(net664),
    .X(_0860_));
 sky130_fd_sc_hd__mux2_1 _1470_ (.A0(net665),
    .A1(\reg_temp[81] ),
    .S(net737),
    .X(_0346_));
 sky130_fd_sc_hd__a221o_1 _1471_ (.A1(net142),
    .A2(net564),
    .B1(net577),
    .B2(\reg_temp[81] ),
    .C1(net928),
    .X(_0861_));
 sky130_fd_sc_hd__mux2_1 _1472_ (.A0(_0861_),
    .A1(\reg_temp[80] ),
    .S(net538),
    .X(_0345_));
 sky130_fd_sc_hd__a221o_1 _1473_ (.A1(net140),
    .A2(net570),
    .B1(net583),
    .B2(\reg_temp[80] ),
    .C1(net826),
    .X(_0862_));
 sky130_fd_sc_hd__mux2_1 _1474_ (.A0(net827),
    .A1(\reg_temp[79] ),
    .S(net538),
    .X(_0344_));
 sky130_fd_sc_hd__a221o_1 _1475_ (.A1(net139),
    .A2(net570),
    .B1(net583),
    .B2(\reg_temp[79] ),
    .C1(net888),
    .X(_0863_));
 sky130_fd_sc_hd__mux2_1 _1476_ (.A0(net889),
    .A1(\reg_temp[78] ),
    .S(net538),
    .X(_0343_));
 sky130_fd_sc_hd__a221o_1 _1477_ (.A1(net138),
    .A2(net569),
    .B1(net582),
    .B2(\reg_temp[78] ),
    .C1(net955),
    .X(_0864_));
 sky130_fd_sc_hd__mux2_1 _1478_ (.A0(net956),
    .A1(\reg_temp[77] ),
    .S(net538),
    .X(_0342_));
 sky130_fd_sc_hd__a221o_1 _1479_ (.A1(net137),
    .A2(net568),
    .B1(net581),
    .B2(\reg_temp[77] ),
    .C1(net1072),
    .X(_0865_));
 sky130_fd_sc_hd__mux2_1 _1480_ (.A0(_0865_),
    .A1(\reg_temp[76] ),
    .S(net538),
    .X(_0341_));
 sky130_fd_sc_hd__a221o_1 _1481_ (.A1(net136),
    .A2(net568),
    .B1(net581),
    .B2(\reg_temp[76] ),
    .C1(net1172),
    .X(_0866_));
 sky130_fd_sc_hd__mux2_1 _1482_ (.A0(net1173),
    .A1(net1433),
    .S(net538),
    .X(_0340_));
 sky130_fd_sc_hd__a221o_1 _1483_ (.A1(net135),
    .A2(net568),
    .B1(net581),
    .B2(\reg_temp[75] ),
    .C1(net1100),
    .X(_0867_));
 sky130_fd_sc_hd__mux2_1 _1484_ (.A0(_0867_),
    .A1(\reg_temp[74] ),
    .S(net538),
    .X(_0339_));
 sky130_fd_sc_hd__a221o_1 _1485_ (.A1(net134),
    .A2(net568),
    .B1(net581),
    .B2(\reg_temp[74] ),
    .C1(net1079),
    .X(_0868_));
 sky130_fd_sc_hd__mux2_1 _1486_ (.A0(net1080),
    .A1(net1567),
    .S(net538),
    .X(_0338_));
 sky130_fd_sc_hd__a221o_1 _1487_ (.A1(net133),
    .A2(net568),
    .B1(net581),
    .B2(\reg_temp[73] ),
    .C1(net1005),
    .X(_0869_));
 sky130_fd_sc_hd__mux2_1 _1488_ (.A0(net1006),
    .A1(\reg_temp[72] ),
    .S(net538),
    .X(_0337_));
 sky130_fd_sc_hd__a221o_1 _1489_ (.A1(net132),
    .A2(net568),
    .B1(net581),
    .B2(\reg_temp[72] ),
    .C1(net1041),
    .X(_0870_));
 sky130_fd_sc_hd__mux2_1 _1490_ (.A0(net1042),
    .A1(\reg_temp[71] ),
    .S(net538),
    .X(_0336_));
 sky130_fd_sc_hd__a221o_1 _1491_ (.A1(net131),
    .A2(net569),
    .B1(net582),
    .B2(\reg_temp[71] ),
    .C1(net1067),
    .X(_0871_));
 sky130_fd_sc_hd__mux2_1 _1492_ (.A0(net1068),
    .A1(\reg_temp[70] ),
    .S(net539),
    .X(_0335_));
 sky130_fd_sc_hd__a221o_1 _1493_ (.A1(net129),
    .A2(net568),
    .B1(net581),
    .B2(\reg_temp[70] ),
    .C1(net1093),
    .X(_0872_));
 sky130_fd_sc_hd__mux2_1 _1494_ (.A0(net1094),
    .A1(\reg_temp[69] ),
    .S(net538),
    .X(_0334_));
 sky130_fd_sc_hd__a221o_1 _1495_ (.A1(net128),
    .A2(net569),
    .B1(net582),
    .B2(\reg_temp[69] ),
    .C1(net1016),
    .X(_0873_));
 sky130_fd_sc_hd__mux2_1 _1496_ (.A0(_0873_),
    .A1(\reg_temp[68] ),
    .S(net538),
    .X(_0333_));
 sky130_fd_sc_hd__a221o_1 _1497_ (.A1(net127),
    .A2(net570),
    .B1(net583),
    .B2(\reg_temp[68] ),
    .C1(net1036),
    .X(_0874_));
 sky130_fd_sc_hd__mux2_1 _1498_ (.A0(net1037),
    .A1(\reg_temp[67] ),
    .S(net538),
    .X(_0332_));
 sky130_fd_sc_hd__a221o_1 _1499_ (.A1(net126),
    .A2(net570),
    .B1(net583),
    .B2(\reg_temp[67] ),
    .C1(net969),
    .X(_0875_));
 sky130_fd_sc_hd__mux2_1 _1500_ (.A0(_0875_),
    .A1(\reg_temp[66] ),
    .S(net538),
    .X(_0331_));
 sky130_fd_sc_hd__a221o_1 _1501_ (.A1(net125),
    .A2(net568),
    .B1(net581),
    .B2(\reg_temp[66] ),
    .C1(net982),
    .X(_0876_));
 sky130_fd_sc_hd__mux2_1 _1502_ (.A0(_0876_),
    .A1(\reg_temp[65] ),
    .S(net538),
    .X(_0330_));
 sky130_fd_sc_hd__a221o_1 _1503_ (.A1(net124),
    .A2(net568),
    .B1(net581),
    .B2(\reg_temp[65] ),
    .C1(net974),
    .X(_0877_));
 sky130_fd_sc_hd__mux2_1 _1504_ (.A0(_0877_),
    .A1(\reg_temp[64] ),
    .S(net538),
    .X(_0329_));
 sky130_fd_sc_hd__a221o_1 _1505_ (.A1(net123),
    .A2(net571),
    .B1(net584),
    .B2(\reg_temp[64] ),
    .C1(net1132),
    .X(_0878_));
 sky130_fd_sc_hd__mux2_1 _1506_ (.A0(net1133),
    .A1(\reg_temp[63] ),
    .S(net539),
    .X(_0328_));
 sky130_fd_sc_hd__a221o_1 _1507_ (.A1(net122),
    .A2(net571),
    .B1(net584),
    .B2(\reg_temp[63] ),
    .C1(net964),
    .X(_0879_));
 sky130_fd_sc_hd__mux2_1 _1508_ (.A0(net965),
    .A1(\reg_temp[62] ),
    .S(net539),
    .X(_0327_));
 sky130_fd_sc_hd__a221o_1 _1509_ (.A1(net121),
    .A2(net571),
    .B1(net584),
    .B2(\reg_temp[62] ),
    .C1(net1030),
    .X(_0880_));
 sky130_fd_sc_hd__mux2_1 _1510_ (.A0(_0880_),
    .A1(net1571),
    .S(net539),
    .X(_0326_));
 sky130_fd_sc_hd__a221o_1 _1511_ (.A1(net120),
    .A2(net571),
    .B1(net584),
    .B2(\reg_temp[61] ),
    .C1(net1157),
    .X(_0881_));
 sky130_fd_sc_hd__mux2_1 _1512_ (.A0(_0881_),
    .A1(\reg_temp[60] ),
    .S(net539),
    .X(_0325_));
 sky130_fd_sc_hd__a221o_1 _1513_ (.A1(net118),
    .A2(net571),
    .B1(net584),
    .B2(\reg_temp[60] ),
    .C1(net1120),
    .X(_0882_));
 sky130_fd_sc_hd__mux2_1 _1514_ (.A0(net1121),
    .A1(\reg_temp[59] ),
    .S(net539),
    .X(_0324_));
 sky130_fd_sc_hd__a221o_1 _1515_ (.A1(net117),
    .A2(net571),
    .B1(net584),
    .B2(\reg_temp[59] ),
    .C1(net1127),
    .X(_0883_));
 sky130_fd_sc_hd__mux2_1 _1516_ (.A0(net1128),
    .A1(\reg_temp[58] ),
    .S(net539),
    .X(_0323_));
 sky130_fd_sc_hd__a221o_1 _1517_ (.A1(net116),
    .A2(net566),
    .B1(net579),
    .B2(\reg_temp[58] ),
    .C1(net997),
    .X(_0884_));
 sky130_fd_sc_hd__mux2_1 _1518_ (.A0(_0884_),
    .A1(net1602),
    .S(net539),
    .X(_0322_));
 sky130_fd_sc_hd__a221o_1 _1519_ (.A1(net115),
    .A2(net571),
    .B1(net584),
    .B2(\reg_temp[57] ),
    .C1(net1107),
    .X(_0885_));
 sky130_fd_sc_hd__mux2_1 _1520_ (.A0(_0885_),
    .A1(\reg_temp[56] ),
    .S(net539),
    .X(_0321_));
 sky130_fd_sc_hd__a221o_1 _1521_ (.A1(net114),
    .A2(net567),
    .B1(net580),
    .B2(\reg_temp[56] ),
    .C1(net1048),
    .X(_0886_));
 sky130_fd_sc_hd__mux2_1 _1522_ (.A0(net1049),
    .A1(\reg_temp[55] ),
    .S(net737),
    .X(_0320_));
 sky130_fd_sc_hd__a221o_1 _1523_ (.A1(net113),
    .A2(net567),
    .B1(net580),
    .B2(\reg_temp[55] ),
    .C1(net1058),
    .X(_0887_));
 sky130_fd_sc_hd__mux2_1 _1524_ (.A0(net1059),
    .A1(\reg_temp[54] ),
    .S(net737),
    .X(_0319_));
 sky130_fd_sc_hd__a221o_1 _1525_ (.A1(net112),
    .A2(net567),
    .B1(net580),
    .B2(\reg_temp[54] ),
    .C1(net1010),
    .X(_0888_));
 sky130_fd_sc_hd__mux2_1 _1526_ (.A0(_0888_),
    .A1(\reg_temp[53] ),
    .S(net737),
    .X(_0318_));
 sky130_fd_sc_hd__a221o_1 _1527_ (.A1(net111),
    .A2(net567),
    .B1(net580),
    .B2(\reg_temp[53] ),
    .C1(net942),
    .X(_0889_));
 sky130_fd_sc_hd__mux2_1 _1528_ (.A0(_0889_),
    .A1(\reg_temp[52] ),
    .S(net737),
    .X(_0317_));
 sky130_fd_sc_hd__a221o_1 _1529_ (.A1(net110),
    .A2(net566),
    .B1(net579),
    .B2(\reg_temp[52] ),
    .C1(net923),
    .X(_0890_));
 sky130_fd_sc_hd__mux2_1 _1530_ (.A0(_0890_),
    .A1(\reg_temp[51] ),
    .S(net770),
    .X(_0316_));
 sky130_fd_sc_hd__a221o_1 _1531_ (.A1(net109),
    .A2(net565),
    .B1(net578),
    .B2(\reg_temp[51] ),
    .C1(net821),
    .X(_0891_));
 sky130_fd_sc_hd__mux2_1 _1532_ (.A0(_0891_),
    .A1(\reg_temp[50] ),
    .S(net737),
    .X(_0315_));
 sky130_fd_sc_hd__a221o_1 _1533_ (.A1(net107),
    .A2(net565),
    .B1(net578),
    .B2(\reg_temp[50] ),
    .C1(net804),
    .X(_0892_));
 sky130_fd_sc_hd__mux2_1 _1534_ (.A0(net805),
    .A1(net1587),
    .S(net737),
    .X(_0314_));
 sky130_fd_sc_hd__a221o_1 _1535_ (.A1(net106),
    .A2(net564),
    .B1(net577),
    .B2(\reg_temp[49] ),
    .C1(net798),
    .X(_0893_));
 sky130_fd_sc_hd__mux2_1 _1536_ (.A0(_0893_),
    .A1(\reg_temp[48] ),
    .S(net737),
    .X(_0313_));
 sky130_fd_sc_hd__a221o_1 _1537_ (.A1(net105),
    .A2(net564),
    .B1(net577),
    .B2(\reg_temp[48] ),
    .C1(net752),
    .X(_0894_));
 sky130_fd_sc_hd__mux2_1 _1538_ (.A0(_0894_),
    .A1(\reg_temp[47] ),
    .S(net737),
    .X(_0312_));
 sky130_fd_sc_hd__a221o_1 _1539_ (.A1(net104),
    .A2(net564),
    .B1(net577),
    .B2(\reg_temp[47] ),
    .C1(net716),
    .X(_0895_));
 sky130_fd_sc_hd__mux2_1 _1540_ (.A0(_0895_),
    .A1(\reg_temp[46] ),
    .S(net737),
    .X(_0311_));
 sky130_fd_sc_hd__a221o_1 _1541_ (.A1(net103),
    .A2(net564),
    .B1(net577),
    .B2(\reg_temp[46] ),
    .C1(net669),
    .X(_0896_));
 sky130_fd_sc_hd__mux2_1 _1542_ (.A0(_0896_),
    .A1(\reg_temp[45] ),
    .S(net737),
    .X(_0310_));
 sky130_fd_sc_hd__a221o_1 _1543_ (.A1(net102),
    .A2(net560),
    .B1(net573),
    .B2(\reg_temp[45] ),
    .C1(net854),
    .X(_0897_));
 sky130_fd_sc_hd__mux2_1 _1544_ (.A0(_0897_),
    .A1(\reg_temp[44] ),
    .S(net737),
    .X(_0309_));
 sky130_fd_sc_hd__a221o_1 _1545_ (.A1(net101),
    .A2(net560),
    .B1(net573),
    .B2(\reg_temp[44] ),
    .C1(net701),
    .X(_0898_));
 sky130_fd_sc_hd__mux2_1 _1546_ (.A0(_0898_),
    .A1(net1454),
    .S(net534),
    .X(_0308_));
 sky130_fd_sc_hd__a221o_1 _1547_ (.A1(net100),
    .A2(net559),
    .B1(net572),
    .B2(\reg_temp[43] ),
    .C1(net729),
    .X(_0899_));
 sky130_fd_sc_hd__mux2_1 _1548_ (.A0(_0899_),
    .A1(\reg_temp[42] ),
    .S(net534),
    .X(_0307_));
 sky130_fd_sc_hd__a221o_1 _1549_ (.A1(net99),
    .A2(net559),
    .B1(net572),
    .B2(\reg_temp[42] ),
    .C1(net840),
    .X(_0900_));
 sky130_fd_sc_hd__mux2_1 _1550_ (.A0(net841),
    .A1(net1646),
    .S(net534),
    .X(_0306_));
 sky130_fd_sc_hd__a221o_1 _1551_ (.A1(net98),
    .A2(net559),
    .B1(net572),
    .B2(\reg_temp[41] ),
    .C1(net848),
    .X(_0901_));
 sky130_fd_sc_hd__mux2_1 _1552_ (.A0(net849),
    .A1(net1648),
    .S(net534),
    .X(_0305_));
 sky130_fd_sc_hd__a221o_1 _1553_ (.A1(net96),
    .A2(net559),
    .B1(net572),
    .B2(\reg_temp[40] ),
    .C1(net911),
    .X(_0902_));
 sky130_fd_sc_hd__mux2_1 _1554_ (.A0(_0902_),
    .A1(net1443),
    .S(net534),
    .X(_0304_));
 sky130_fd_sc_hd__a221o_1 _1555_ (.A1(net95),
    .A2(net559),
    .B1(net572),
    .B2(\reg_temp[39] ),
    .C1(net884),
    .X(_0903_));
 sky130_fd_sc_hd__mux2_1 _1556_ (.A0(_0903_),
    .A1(net1450),
    .S(net737),
    .X(_0303_));
 sky130_fd_sc_hd__a221o_1 _1557_ (.A1(net94),
    .A2(net561),
    .B1(net574),
    .B2(\reg_temp[38] ),
    .C1(net993),
    .X(_0904_));
 sky130_fd_sc_hd__mux2_1 _1558_ (.A0(_0904_),
    .A1(\reg_temp[37] ),
    .S(net738),
    .X(_0302_));
 sky130_fd_sc_hd__a221o_1 _1559_ (.A1(net93),
    .A2(net561),
    .B1(net574),
    .B2(\reg_temp[37] ),
    .C1(net1001),
    .X(_0905_));
 sky130_fd_sc_hd__mux2_1 _1560_ (.A0(net1002),
    .A1(net1607),
    .S(net738),
    .X(_0301_));
 sky130_fd_sc_hd__a221o_1 _1561_ (.A1(net92),
    .A2(net561),
    .B1(net574),
    .B2(\reg_temp[36] ),
    .C1(net1026),
    .X(_0906_));
 sky130_fd_sc_hd__mux2_1 _1562_ (.A0(net1027),
    .A1(net1644),
    .S(net738),
    .X(_0300_));
 sky130_fd_sc_hd__a221o_1 _1563_ (.A1(net91),
    .A2(net563),
    .B1(net576),
    .B2(\reg_temp[35] ),
    .C1(net793),
    .X(_0907_));
 sky130_fd_sc_hd__mux2_1 _1564_ (.A0(net794),
    .A1(net1597),
    .S(net738),
    .X(_0299_));
 sky130_fd_sc_hd__a221o_1 _1565_ (.A1(net90),
    .A2(net563),
    .B1(net576),
    .B2(\reg_temp[34] ),
    .C1(net763),
    .X(_0908_));
 sky130_fd_sc_hd__mux2_1 _1566_ (.A0(_0908_),
    .A1(net1590),
    .S(net738),
    .X(_0298_));
 sky130_fd_sc_hd__a221o_1 _1567_ (.A1(net89),
    .A2(net563),
    .B1(net576),
    .B2(\reg_temp[33] ),
    .C1(net1063),
    .X(_0909_));
 sky130_fd_sc_hd__mux2_1 _1568_ (.A0(net1064),
    .A1(net1578),
    .S(net738),
    .X(_0297_));
 sky130_fd_sc_hd__a221o_1 _1569_ (.A1(net88),
    .A2(net563),
    .B1(net576),
    .B2(\reg_temp[32] ),
    .C1(net901),
    .X(_0910_));
 sky130_fd_sc_hd__mux2_1 _1570_ (.A0(net902),
    .A1(net1594),
    .S(net738),
    .X(_0296_));
 sky130_fd_sc_hd__a221o_1 _1571_ (.A1(net87),
    .A2(net561),
    .B1(net574),
    .B2(\reg_temp[31] ),
    .C1(net933),
    .X(_0911_));
 sky130_fd_sc_hd__mux2_1 _1572_ (.A0(_0911_),
    .A1(net1586),
    .S(net738),
    .X(_0295_));
 sky130_fd_sc_hd__a221o_1 _1573_ (.A1(net85),
    .A2(net562),
    .B1(net575),
    .B2(\reg_temp[30] ),
    .C1(net947),
    .X(_0912_));
 sky130_fd_sc_hd__mux2_1 _1574_ (.A0(net948),
    .A1(net1639),
    .S(net738),
    .X(_0294_));
 sky130_fd_sc_hd__a221o_1 _1575_ (.A1(net84),
    .A2(net562),
    .B1(net575),
    .B2(\reg_temp[29] ),
    .C1(net880),
    .X(_0913_));
 sky130_fd_sc_hd__mux2_1 _1576_ (.A0(net881),
    .A1(net1619),
    .S(net535),
    .X(_0293_));
 sky130_fd_sc_hd__a221o_1 _1577_ (.A1(net83),
    .A2(net562),
    .B1(net575),
    .B2(\reg_temp[28] ),
    .C1(net894),
    .X(_0914_));
 sky130_fd_sc_hd__mux2_1 _1578_ (.A0(net895),
    .A1(net1613),
    .S(net535),
    .X(_0292_));
 sky130_fd_sc_hd__a221o_1 _1579_ (.A1(net82),
    .A2(net562),
    .B1(net575),
    .B2(\reg_temp[27] ),
    .C1(net905),
    .X(_0915_));
 sky130_fd_sc_hd__mux2_1 _1580_ (.A0(_0915_),
    .A1(net1595),
    .S(net535),
    .X(_0291_));
 sky130_fd_sc_hd__a221o_1 _1581_ (.A1(net81),
    .A2(net561),
    .B1(net574),
    .B2(\reg_temp[26] ),
    .C1(net865),
    .X(_0916_));
 sky130_fd_sc_hd__mux2_1 _1582_ (.A0(net866),
    .A1(net1626),
    .S(net535),
    .X(_0290_));
 sky130_fd_sc_hd__a221o_1 _1583_ (.A1(net80),
    .A2(net561),
    .B1(net574),
    .B2(\reg_temp[25] ),
    .C1(net784),
    .X(_0917_));
 sky130_fd_sc_hd__mux2_1 _1584_ (.A0(_0917_),
    .A1(net1584),
    .S(net535),
    .X(_0289_));
 sky130_fd_sc_hd__a221o_1 _1585_ (.A1(net79),
    .A2(net561),
    .B1(net574),
    .B2(\reg_temp[24] ),
    .C1(net1193),
    .X(_0918_));
 sky130_fd_sc_hd__mux2_1 _1586_ (.A0(_0918_),
    .A1(net1647),
    .S(net534),
    .X(_0288_));
 sky130_fd_sc_hd__a221o_1 _1587_ (.A1(net78),
    .A2(net562),
    .B1(net575),
    .B2(\reg_temp[23] ),
    .C1(net1182),
    .X(_0919_));
 sky130_fd_sc_hd__mux2_1 _1588_ (.A0(net1183),
    .A1(net1638),
    .S(net535),
    .X(_0287_));
 sky130_fd_sc_hd__a221o_1 _1589_ (.A1(net77),
    .A2(net561),
    .B1(net575),
    .B2(\reg_temp[22] ),
    .C1(net1186),
    .X(_0920_));
 sky130_fd_sc_hd__mux2_1 _1590_ (.A0(net1187),
    .A1(net1630),
    .S(net738),
    .X(_0286_));
 sky130_fd_sc_hd__a221o_1 _1591_ (.A1(net76),
    .A2(net561),
    .B1(net574),
    .B2(\reg_temp[21] ),
    .C1(net1178),
    .X(_0921_));
 sky130_fd_sc_hd__mux2_1 _1592_ (.A0(_0921_),
    .A1(net1637),
    .S(net535),
    .X(_0285_));
 sky130_fd_sc_hd__a221o_1 _1593_ (.A1(net74),
    .A2(net562),
    .B1(net574),
    .B2(\reg_temp[20] ),
    .C1(_0806_),
    .X(_0922_));
 sky130_fd_sc_hd__mux2_1 _1594_ (.A0(_0922_),
    .A1(net1621),
    .S(net535),
    .X(_0284_));
 sky130_fd_sc_hd__a221o_1 _1595_ (.A1(net73),
    .A2(net562),
    .B1(net574),
    .B2(\reg_temp[19] ),
    .C1(_0808_),
    .X(_0923_));
 sky130_fd_sc_hd__mux2_1 _1596_ (.A0(_0923_),
    .A1(net1620),
    .S(net535),
    .X(_0283_));
 sky130_fd_sc_hd__a221o_1 _1597_ (.A1(net72),
    .A2(net562),
    .B1(net575),
    .B2(\reg_temp[18] ),
    .C1(_0810_),
    .X(_0924_));
 sky130_fd_sc_hd__mux2_1 _1598_ (.A0(_0924_),
    .A1(net1642),
    .S(net535),
    .X(_0282_));
 sky130_fd_sc_hd__a221o_1 _1599_ (.A1(net71),
    .A2(net562),
    .B1(net575),
    .B2(\reg_temp[17] ),
    .C1(net1169),
    .X(_0925_));
 sky130_fd_sc_hd__mux2_1 _1600_ (.A0(_0925_),
    .A1(\reg_temp[16] ),
    .S(net535),
    .X(_0281_));
 sky130_fd_sc_hd__a221o_1 _1601_ (.A1(net67),
    .A2(net561),
    .B1(net574),
    .B2(\reg_temp[16] ),
    .C1(net789),
    .X(_0926_));
 sky130_fd_sc_hd__mux2_1 _1602_ (.A0(_0926_),
    .A1(net1599),
    .S(net535),
    .X(_0280_));
 sky130_fd_sc_hd__a221o_1 _1603_ (.A1(net56),
    .A2(net561),
    .B1(net574),
    .B2(\reg_temp[15] ),
    .C1(net742),
    .X(_0927_));
 sky130_fd_sc_hd__mux2_1 _1604_ (.A0(_0927_),
    .A1(\reg_temp[14] ),
    .S(net535),
    .X(_0279_));
 sky130_fd_sc_hd__a221o_1 _1605_ (.A1(net45),
    .A2(net561),
    .B1(net574),
    .B2(\reg_temp[14] ),
    .C1(net876),
    .X(_0928_));
 sky130_fd_sc_hd__mux2_1 _1606_ (.A0(net877),
    .A1(net1629),
    .S(net534),
    .X(_0278_));
 sky130_fd_sc_hd__a221o_1 _1607_ (.A1(net34),
    .A2(net561),
    .B1(net574),
    .B2(\reg_temp[13] ),
    .C1(net860),
    .X(_0929_));
 sky130_fd_sc_hd__mux2_1 _1608_ (.A0(net861),
    .A1(net1589),
    .S(net534),
    .X(_0277_));
 sky130_fd_sc_hd__a221o_1 _1609_ (.A1(net23),
    .A2(net559),
    .B1(net572),
    .B2(\reg_temp[12] ),
    .C1(net813),
    .X(_0930_));
 sky130_fd_sc_hd__mux2_1 _1610_ (.A0(net814),
    .A1(\reg_temp[11] ),
    .S(net737),
    .X(_0276_));
 sky130_fd_sc_hd__a221o_1 _1611_ (.A1(net12),
    .A2(net559),
    .B1(net572),
    .B2(\reg_temp[11] ),
    .C1(net711),
    .X(_0931_));
 sky130_fd_sc_hd__mux2_1 _1612_ (.A0(net712),
    .A1(\reg_temp[10] ),
    .S(net534),
    .X(_0275_));
 sky130_fd_sc_hd__a221o_1 _1613_ (.A1(net163),
    .A2(net559),
    .B1(net572),
    .B2(\reg_temp[10] ),
    .C1(net758),
    .X(_0932_));
 sky130_fd_sc_hd__mux2_1 _1614_ (.A0(net759),
    .A1(\reg_temp[9] ),
    .S(net534),
    .X(_0274_));
 sky130_fd_sc_hd__a221o_1 _1615_ (.A1(net152),
    .A2(net561),
    .B1(net572),
    .B2(\reg_temp[9] ),
    .C1(net844),
    .X(_0933_));
 sky130_fd_sc_hd__mux2_1 _1616_ (.A0(net845),
    .A1(net1650),
    .S(net534),
    .X(_0273_));
 sky130_fd_sc_hd__a221o_1 _1617_ (.A1(net141),
    .A2(net562),
    .B1(net575),
    .B2(\reg_temp[8] ),
    .C1(net774),
    .X(_0934_));
 sky130_fd_sc_hd__mux2_1 _1618_ (.A0(_0934_),
    .A1(\reg_temp[7] ),
    .S(net535),
    .X(_0272_));
 sky130_fd_sc_hd__a221o_1 _1619_ (.A1(net130),
    .A2(net562),
    .B1(net575),
    .B2(\reg_temp[7] ),
    .C1(net721),
    .X(_0935_));
 sky130_fd_sc_hd__mux2_1 _1620_ (.A0(_0935_),
    .A1(\reg_temp[6] ),
    .S(net535),
    .X(_0271_));
 sky130_fd_sc_hd__a221o_1 _1621_ (.A1(net119),
    .A2(net561),
    .B1(net574),
    .B2(\reg_temp[6] ),
    .C1(net725),
    .X(_0936_));
 sky130_fd_sc_hd__mux2_1 _1622_ (.A0(_0936_),
    .A1(net1615),
    .S(net535),
    .X(_0270_));
 sky130_fd_sc_hd__a221o_1 _1623_ (.A1(net108),
    .A2(net561),
    .B1(net574),
    .B2(\reg_temp[5] ),
    .C1(net938),
    .X(_0937_));
 sky130_fd_sc_hd__mux2_1 _1624_ (.A0(_0937_),
    .A1(net1608),
    .S(net534),
    .X(_0269_));
 sky130_fd_sc_hd__a221o_1 _1625_ (.A1(net97),
    .A2(net559),
    .B1(net572),
    .B2(\reg_temp[4] ),
    .C1(net833),
    .X(_0938_));
 sky130_fd_sc_hd__mux2_1 _1626_ (.A0(net834),
    .A1(net1622),
    .S(net534),
    .X(_0268_));
 sky130_fd_sc_hd__a221o_1 _1627_ (.A1(net86),
    .A2(net559),
    .B1(net572),
    .B2(\reg_temp[3] ),
    .C1(net674),
    .X(_0939_));
 sky130_fd_sc_hd__mux2_1 _1628_ (.A0(net675),
    .A1(\reg_temp[2] ),
    .S(net534),
    .X(_0267_));
 sky130_fd_sc_hd__a221o_1 _1629_ (.A1(net75),
    .A2(net559),
    .B1(net572),
    .B2(\reg_temp[2] ),
    .C1(net688),
    .X(_0940_));
 sky130_fd_sc_hd__mux2_1 _1630_ (.A0(net689),
    .A1(\reg_temp[1] ),
    .S(net534),
    .X(_0266_));
 sky130_fd_sc_hd__a221o_1 _1631_ (.A1(net1),
    .A2(net559),
    .B1(net572),
    .B2(\reg_temp[1] ),
    .C1(net706),
    .X(_0941_));
 sky130_fd_sc_hd__mux2_1 _1632_ (.A0(net707),
    .A1(\reg_temp[0] ),
    .S(net534),
    .X(_0265_));
 sky130_fd_sc_hd__or4b_2 _1633_ (.A(net174),
    .B(net173),
    .C(_0573_),
    .D_N(_0591_),
    .X(_0942_));
 sky130_fd_sc_hd__nand2_1 _1634_ (.A(net176),
    .B(net177),
    .Y(_0943_));
 sky130_fd_sc_hd__or4_1 _1635_ (.A(net179),
    .B(net178),
    .C(net572),
    .D(_0943_),
    .X(_0944_));
 sky130_fd_sc_hd__nor2_1 _1636_ (.A(_0942_),
    .B(_0944_),
    .Y(_0001_));
 sky130_fd_sc_hd__nor2_1 _1637_ (.A(net261),
    .B(net559),
    .Y(_0002_));
 sky130_fd_sc_hd__or3_1 _1638_ (.A(\current_state[0] ),
    .B(\current_state[1] ),
    .C(net515),
    .X(_0945_));
 sky130_fd_sc_hd__o21a_1 _1639_ (.A1(net591),
    .A2(_0002_),
    .B1(_0945_),
    .X(\next_state[0] ));
 sky130_fd_sc_hd__a221o_1 _1640_ (.A1(enable_proc),
    .A2(_0523_),
    .B1(net559),
    .B2(_0522_),
    .C1(net572),
    .X(\next_state[1] ));
 sky130_fd_sc_hd__nor2_1 _1641_ (.A(net441),
    .B(_0524_),
    .Y(_0946_));
 sky130_fd_sc_hd__and2_2 _1642_ (.A(\reg_temp[0] ),
    .B(net540),
    .X(net263));
 sky130_fd_sc_hd__and2_1 _1643_ (.A(\reg_temp[1] ),
    .B(net540),
    .X(net337));
 sky130_fd_sc_hd__and2_1 _1644_ (.A(\reg_temp[2] ),
    .B(net540),
    .X(net348));
 sky130_fd_sc_hd__and2_1 _1645_ (.A(\reg_temp[3] ),
    .B(net540),
    .X(net359));
 sky130_fd_sc_hd__and2_1 _1646_ (.A(\reg_temp[4] ),
    .B(net540),
    .X(net370));
 sky130_fd_sc_hd__and2_1 _1647_ (.A(\reg_temp[5] ),
    .B(net542),
    .X(net381));
 sky130_fd_sc_hd__and2_1 _1648_ (.A(\reg_temp[6] ),
    .B(net541),
    .X(net392));
 sky130_fd_sc_hd__and2_1 _1649_ (.A(\reg_temp[7] ),
    .B(net541),
    .X(net403));
 sky130_fd_sc_hd__and2_1 _1650_ (.A(\reg_temp[8] ),
    .B(net541),
    .X(net414));
 sky130_fd_sc_hd__and2_1 _1651_ (.A(\reg_temp[9] ),
    .B(net540),
    .X(net425));
 sky130_fd_sc_hd__and2_1 _1652_ (.A(\reg_temp[10] ),
    .B(net540),
    .X(net274));
 sky130_fd_sc_hd__and2_1 _1653_ (.A(\reg_temp[11] ),
    .B(net540),
    .X(net285));
 sky130_fd_sc_hd__and2_1 _1654_ (.A(\reg_temp[12] ),
    .B(net540),
    .X(net296));
 sky130_fd_sc_hd__and2_1 _1655_ (.A(\reg_temp[13] ),
    .B(net540),
    .X(net307));
 sky130_fd_sc_hd__and2_1 _1656_ (.A(\reg_temp[14] ),
    .B(net542),
    .X(net318));
 sky130_fd_sc_hd__and2_1 _1657_ (.A(\reg_temp[15] ),
    .B(net542),
    .X(net329));
 sky130_fd_sc_hd__and2_1 _1658_ (.A(\reg_temp[16] ),
    .B(net542),
    .X(net333));
 sky130_fd_sc_hd__and2_1 _1659_ (.A(\reg_temp[17] ),
    .B(net541),
    .X(net334));
 sky130_fd_sc_hd__and2_1 _1660_ (.A(\reg_temp[18] ),
    .B(net541),
    .X(net335));
 sky130_fd_sc_hd__and2_1 _1661_ (.A(\reg_temp[19] ),
    .B(net541),
    .X(net336));
 sky130_fd_sc_hd__and2_1 _1662_ (.A(\reg_temp[20] ),
    .B(net542),
    .X(net338));
 sky130_fd_sc_hd__and2_1 _1663_ (.A(\reg_temp[21] ),
    .B(net542),
    .X(net339));
 sky130_fd_sc_hd__and2_1 _1664_ (.A(\reg_temp[22] ),
    .B(net542),
    .X(net340));
 sky130_fd_sc_hd__and2_1 _1665_ (.A(\reg_temp[23] ),
    .B(net542),
    .X(net341));
 sky130_fd_sc_hd__and2_1 _1666_ (.A(\reg_temp[24] ),
    .B(net542),
    .X(net342));
 sky130_fd_sc_hd__and2_1 _1667_ (.A(\reg_temp[25] ),
    .B(net542),
    .X(net343));
 sky130_fd_sc_hd__and2_1 _1668_ (.A(\reg_temp[26] ),
    .B(net541),
    .X(net344));
 sky130_fd_sc_hd__and2_1 _1669_ (.A(\reg_temp[27] ),
    .B(net541),
    .X(net345));
 sky130_fd_sc_hd__and2_1 _1670_ (.A(\reg_temp[28] ),
    .B(net541),
    .X(net346));
 sky130_fd_sc_hd__and2_1 _1671_ (.A(\reg_temp[29] ),
    .B(net541),
    .X(net347));
 sky130_fd_sc_hd__and2_1 _1672_ (.A(\reg_temp[30] ),
    .B(net541),
    .X(net349));
 sky130_fd_sc_hd__and2_1 _1673_ (.A(\reg_temp[31] ),
    .B(net541),
    .X(net350));
 sky130_fd_sc_hd__and2_1 _1674_ (.A(\reg_temp[32] ),
    .B(net541),
    .X(net351));
 sky130_fd_sc_hd__and2_1 _1675_ (.A(\reg_temp[33] ),
    .B(net541),
    .X(net352));
 sky130_fd_sc_hd__and2_1 _1676_ (.A(\reg_temp[34] ),
    .B(net541),
    .X(net353));
 sky130_fd_sc_hd__and2_1 _1677_ (.A(\reg_temp[35] ),
    .B(net541),
    .X(net354));
 sky130_fd_sc_hd__and2_1 _1678_ (.A(\reg_temp[36] ),
    .B(net542),
    .X(net355));
 sky130_fd_sc_hd__and2_1 _1679_ (.A(\reg_temp[37] ),
    .B(net542),
    .X(net356));
 sky130_fd_sc_hd__and2_1 _1680_ (.A(\reg_temp[38] ),
    .B(net542),
    .X(net357));
 sky130_fd_sc_hd__and2_1 _1681_ (.A(\reg_temp[39] ),
    .B(net540),
    .X(net358));
 sky130_fd_sc_hd__and2_1 _1682_ (.A(\reg_temp[40] ),
    .B(net543),
    .X(net360));
 sky130_fd_sc_hd__and2_2 _1683_ (.A(\reg_temp[41] ),
    .B(net540),
    .X(net361));
 sky130_fd_sc_hd__and2_1 _1684_ (.A(\reg_temp[42] ),
    .B(net540),
    .X(net362));
 sky130_fd_sc_hd__and2_2 _1685_ (.A(\reg_temp[43] ),
    .B(net540),
    .X(net363));
 sky130_fd_sc_hd__and2_1 _1686_ (.A(\reg_temp[44] ),
    .B(net540),
    .X(net364));
 sky130_fd_sc_hd__and2_2 _1687_ (.A(\reg_temp[45] ),
    .B(net544),
    .X(net365));
 sky130_fd_sc_hd__and2_1 _1688_ (.A(\reg_temp[46] ),
    .B(net544),
    .X(net366));
 sky130_fd_sc_hd__and2_1 _1689_ (.A(\reg_temp[47] ),
    .B(net544),
    .X(net367));
 sky130_fd_sc_hd__and2_1 _1690_ (.A(\reg_temp[48] ),
    .B(net544),
    .X(net368));
 sky130_fd_sc_hd__and2_1 _1691_ (.A(\reg_temp[49] ),
    .B(net544),
    .X(net369));
 sky130_fd_sc_hd__and2_1 _1692_ (.A(\reg_temp[50] ),
    .B(net543),
    .X(net371));
 sky130_fd_sc_hd__and2_1 _1693_ (.A(\reg_temp[51] ),
    .B(net543),
    .X(net372));
 sky130_fd_sc_hd__and2_1 _1694_ (.A(\reg_temp[52] ),
    .B(net543),
    .X(net373));
 sky130_fd_sc_hd__and2_1 _1695_ (.A(\reg_temp[53] ),
    .B(net543),
    .X(net374));
 sky130_fd_sc_hd__and2_1 _1696_ (.A(\reg_temp[54] ),
    .B(net543),
    .X(net375));
 sky130_fd_sc_hd__and2_1 _1697_ (.A(\reg_temp[55] ),
    .B(net543),
    .X(net376));
 sky130_fd_sc_hd__and2_1 _1698_ (.A(\reg_temp[56] ),
    .B(net543),
    .X(net377));
 sky130_fd_sc_hd__and2_1 _1699_ (.A(\reg_temp[57] ),
    .B(net543),
    .X(net378));
 sky130_fd_sc_hd__and2_1 _1700_ (.A(\reg_temp[58] ),
    .B(net543),
    .X(net379));
 sky130_fd_sc_hd__and2_1 _1701_ (.A(\reg_temp[59] ),
    .B(net543),
    .X(net380));
 sky130_fd_sc_hd__and2_1 _1702_ (.A(\reg_temp[60] ),
    .B(net543),
    .X(net382));
 sky130_fd_sc_hd__and2_1 _1703_ (.A(\reg_temp[61] ),
    .B(net543),
    .X(net383));
 sky130_fd_sc_hd__and2_1 _1704_ (.A(\reg_temp[62] ),
    .B(net543),
    .X(net384));
 sky130_fd_sc_hd__and2_1 _1705_ (.A(\reg_temp[63] ),
    .B(net544),
    .X(net385));
 sky130_fd_sc_hd__and2_1 _1706_ (.A(\reg_temp[64] ),
    .B(net543),
    .X(net386));
 sky130_fd_sc_hd__and2_1 _1707_ (.A(\reg_temp[65] ),
    .B(net548),
    .X(net387));
 sky130_fd_sc_hd__and2_1 _1708_ (.A(\reg_temp[66] ),
    .B(net546),
    .X(net388));
 sky130_fd_sc_hd__and2_1 _1709_ (.A(\reg_temp[67] ),
    .B(net546),
    .X(net389));
 sky130_fd_sc_hd__and2_2 _1710_ (.A(\reg_temp[68] ),
    .B(net545),
    .X(net390));
 sky130_fd_sc_hd__and2_2 _1711_ (.A(\reg_temp[69] ),
    .B(net545),
    .X(net391));
 sky130_fd_sc_hd__and2_1 _1712_ (.A(\reg_temp[70] ),
    .B(net550),
    .X(net393));
 sky130_fd_sc_hd__and2_1 _1713_ (.A(\reg_temp[71] ),
    .B(net547),
    .X(net394));
 sky130_fd_sc_hd__and2_1 _1714_ (.A(\reg_temp[72] ),
    .B(net547),
    .X(net395));
 sky130_fd_sc_hd__and2_1 _1715_ (.A(\reg_temp[73] ),
    .B(net543),
    .X(net396));
 sky130_fd_sc_hd__and2_1 _1716_ (.A(\reg_temp[74] ),
    .B(net549),
    .X(net397));
 sky130_fd_sc_hd__and2_1 _1717_ (.A(\reg_temp[75] ),
    .B(net549),
    .X(net398));
 sky130_fd_sc_hd__and2_1 _1718_ (.A(\reg_temp[76] ),
    .B(net548),
    .X(net399));
 sky130_fd_sc_hd__and2_1 _1719_ (.A(\reg_temp[77] ),
    .B(net547),
    .X(net400));
 sky130_fd_sc_hd__and2_1 _1720_ (.A(\reg_temp[78] ),
    .B(net550),
    .X(net401));
 sky130_fd_sc_hd__and2_2 _1721_ (.A(\reg_temp[79] ),
    .B(net545),
    .X(net402));
 sky130_fd_sc_hd__and2_1 _1722_ (.A(\reg_temp[80] ),
    .B(net545),
    .X(net404));
 sky130_fd_sc_hd__and2_2 _1723_ (.A(\reg_temp[81] ),
    .B(net546),
    .X(net405));
 sky130_fd_sc_hd__and2_2 _1724_ (.A(\reg_temp[82] ),
    .B(net544),
    .X(net406));
 sky130_fd_sc_hd__and2_2 _1725_ (.A(\reg_temp[83] ),
    .B(net540),
    .X(net407));
 sky130_fd_sc_hd__and2_1 _1726_ (.A(\reg_temp[84] ),
    .B(net546),
    .X(net408));
 sky130_fd_sc_hd__and2_1 _1727_ (.A(\reg_temp[85] ),
    .B(net546),
    .X(net409));
 sky130_fd_sc_hd__and2_1 _1728_ (.A(\reg_temp[86] ),
    .B(net548),
    .X(net410));
 sky130_fd_sc_hd__and2_1 _1729_ (.A(\reg_temp[87] ),
    .B(net548),
    .X(net411));
 sky130_fd_sc_hd__and2_1 _1730_ (.A(\reg_temp[88] ),
    .B(net548),
    .X(net412));
 sky130_fd_sc_hd__and2_1 _1731_ (.A(\reg_temp[89] ),
    .B(net547),
    .X(net413));
 sky130_fd_sc_hd__and2_1 _1732_ (.A(\reg_temp[90] ),
    .B(net547),
    .X(net415));
 sky130_fd_sc_hd__and2_2 _1733_ (.A(\reg_temp[91] ),
    .B(net546),
    .X(net416));
 sky130_fd_sc_hd__and2_1 _1734_ (.A(\reg_temp[92] ),
    .B(net546),
    .X(net417));
 sky130_fd_sc_hd__and2_1 _1735_ (.A(\reg_temp[93] ),
    .B(net546),
    .X(net418));
 sky130_fd_sc_hd__and2_1 _1736_ (.A(\reg_temp[94] ),
    .B(net546),
    .X(net419));
 sky130_fd_sc_hd__and2_2 _1737_ (.A(\reg_temp[95] ),
    .B(net546),
    .X(net420));
 sky130_fd_sc_hd__and2_1 _1738_ (.A(\reg_temp[96] ),
    .B(net548),
    .X(net421));
 sky130_fd_sc_hd__and2_1 _1739_ (.A(\reg_temp[97] ),
    .B(net548),
    .X(net422));
 sky130_fd_sc_hd__and2_1 _1740_ (.A(\reg_temp[98] ),
    .B(net548),
    .X(net423));
 sky130_fd_sc_hd__and2_1 _1741_ (.A(\reg_temp[99] ),
    .B(net547),
    .X(net424));
 sky130_fd_sc_hd__and2_1 _1742_ (.A(\reg_temp[100] ),
    .B(net547),
    .X(net264));
 sky130_fd_sc_hd__and2_1 _1743_ (.A(\reg_temp[101] ),
    .B(net547),
    .X(net265));
 sky130_fd_sc_hd__and2_1 _1744_ (.A(\reg_temp[102] ),
    .B(net547),
    .X(net266));
 sky130_fd_sc_hd__and2_1 _1745_ (.A(\reg_temp[103] ),
    .B(net547),
    .X(net267));
 sky130_fd_sc_hd__and2_1 _1746_ (.A(\reg_temp[104] ),
    .B(net547),
    .X(net268));
 sky130_fd_sc_hd__and2_1 _1747_ (.A(\reg_temp[105] ),
    .B(net547),
    .X(net269));
 sky130_fd_sc_hd__and2_1 _1748_ (.A(\reg_temp[106] ),
    .B(net548),
    .X(net270));
 sky130_fd_sc_hd__and2_1 _1749_ (.A(\reg_temp[107] ),
    .B(net548),
    .X(net271));
 sky130_fd_sc_hd__and2_1 _1750_ (.A(\reg_temp[108] ),
    .B(net548),
    .X(net272));
 sky130_fd_sc_hd__and2_1 _1751_ (.A(\reg_temp[109] ),
    .B(net551),
    .X(net273));
 sky130_fd_sc_hd__and2_1 _1752_ (.A(\reg_temp[110] ),
    .B(net548),
    .X(net275));
 sky130_fd_sc_hd__and2_1 _1753_ (.A(\reg_temp[111] ),
    .B(net547),
    .X(net276));
 sky130_fd_sc_hd__and2_1 _1754_ (.A(\reg_temp[112] ),
    .B(net547),
    .X(net277));
 sky130_fd_sc_hd__and2_1 _1755_ (.A(\reg_temp[113] ),
    .B(net547),
    .X(net278));
 sky130_fd_sc_hd__and2_1 _1756_ (.A(\reg_temp[114] ),
    .B(net547),
    .X(net279));
 sky130_fd_sc_hd__and2_1 _1757_ (.A(\reg_temp[115] ),
    .B(net551),
    .X(net280));
 sky130_fd_sc_hd__and2_1 _1758_ (.A(\reg_temp[116] ),
    .B(net548),
    .X(net281));
 sky130_fd_sc_hd__and2_1 _1759_ (.A(\reg_temp[117] ),
    .B(net551),
    .X(net282));
 sky130_fd_sc_hd__and2_1 _1760_ (.A(\reg_temp[118] ),
    .B(net548),
    .X(net283));
 sky130_fd_sc_hd__and2_1 _1761_ (.A(\reg_temp[119] ),
    .B(net548),
    .X(net284));
 sky130_fd_sc_hd__and2_1 _1762_ (.A(\reg_temp[120] ),
    .B(net546),
    .X(net286));
 sky130_fd_sc_hd__and2_1 _1763_ (.A(\reg_temp[121] ),
    .B(net546),
    .X(net287));
 sky130_fd_sc_hd__and2_2 _1764_ (.A(\reg_temp[122] ),
    .B(net546),
    .X(net288));
 sky130_fd_sc_hd__and2_1 _1765_ (.A(\reg_temp[123] ),
    .B(net546),
    .X(net289));
 sky130_fd_sc_hd__and2_1 _1766_ (.A(\reg_temp[124] ),
    .B(net546),
    .X(net290));
 sky130_fd_sc_hd__and2_2 _1767_ (.A(\reg_temp[125] ),
    .B(net545),
    .X(net291));
 sky130_fd_sc_hd__and2_2 _1768_ (.A(\reg_temp[126] ),
    .B(net545),
    .X(net292));
 sky130_fd_sc_hd__and2_1 _1769_ (.A(\reg_temp[127] ),
    .B(net545),
    .X(net293));
 sky130_fd_sc_hd__and2_1 _1770_ (.A(\reg_temp[128] ),
    .B(net545),
    .X(net294));
 sky130_fd_sc_hd__and2_1 _1771_ (.A(\reg_temp[129] ),
    .B(net545),
    .X(net295));
 sky130_fd_sc_hd__and2_1 _1772_ (.A(\reg_temp[130] ),
    .B(net551),
    .X(net297));
 sky130_fd_sc_hd__and2_1 _1773_ (.A(\reg_temp[131] ),
    .B(net545),
    .X(net298));
 sky130_fd_sc_hd__and2_1 _1774_ (.A(\reg_temp[132] ),
    .B(net545),
    .X(net299));
 sky130_fd_sc_hd__and2_1 _1775_ (.A(\reg_temp[133] ),
    .B(net550),
    .X(net300));
 sky130_fd_sc_hd__and2_1 _1776_ (.A(\reg_temp[134] ),
    .B(net550),
    .X(net301));
 sky130_fd_sc_hd__and2_1 _1777_ (.A(\reg_temp[135] ),
    .B(net549),
    .X(net302));
 sky130_fd_sc_hd__and2_1 _1778_ (.A(\reg_temp[136] ),
    .B(net549),
    .X(net303));
 sky130_fd_sc_hd__and2_1 _1779_ (.A(\reg_temp[137] ),
    .B(net549),
    .X(net304));
 sky130_fd_sc_hd__and2_1 _1780_ (.A(\reg_temp[138] ),
    .B(net549),
    .X(net305));
 sky130_fd_sc_hd__and2_1 _1781_ (.A(\reg_temp[139] ),
    .B(net549),
    .X(net306));
 sky130_fd_sc_hd__and2_1 _1782_ (.A(\reg_temp[140] ),
    .B(net550),
    .X(net308));
 sky130_fd_sc_hd__and2_1 _1783_ (.A(\reg_temp[141] ),
    .B(net549),
    .X(net309));
 sky130_fd_sc_hd__and2_1 _1784_ (.A(\reg_temp[142] ),
    .B(net549),
    .X(net310));
 sky130_fd_sc_hd__and2_1 _1785_ (.A(\reg_temp[143] ),
    .B(net549),
    .X(net311));
 sky130_fd_sc_hd__and2_1 _1786_ (.A(\reg_temp[144] ),
    .B(net549),
    .X(net312));
 sky130_fd_sc_hd__and2_1 _1787_ (.A(\reg_temp[145] ),
    .B(net549),
    .X(net313));
 sky130_fd_sc_hd__and2_1 _1788_ (.A(\reg_temp[146] ),
    .B(net550),
    .X(net314));
 sky130_fd_sc_hd__and2_1 _1789_ (.A(\reg_temp[147] ),
    .B(net550),
    .X(net315));
 sky130_fd_sc_hd__and2_1 _1790_ (.A(\reg_temp[148] ),
    .B(net545),
    .X(net316));
 sky130_fd_sc_hd__and2_1 _1791_ (.A(\reg_temp[149] ),
    .B(net545),
    .X(net317));
 sky130_fd_sc_hd__and2_1 _1792_ (.A(\reg_temp[150] ),
    .B(net551),
    .X(net319));
 sky130_fd_sc_hd__and2_1 _1793_ (.A(\reg_temp[151] ),
    .B(net545),
    .X(net320));
 sky130_fd_sc_hd__and2_1 _1794_ (.A(\reg_temp[152] ),
    .B(net550),
    .X(net321));
 sky130_fd_sc_hd__and2_1 _1795_ (.A(\reg_temp[153] ),
    .B(net549),
    .X(net322));
 sky130_fd_sc_hd__and2_1 _1796_ (.A(\reg_temp[154] ),
    .B(net549),
    .X(net323));
 sky130_fd_sc_hd__and2_1 _1797_ (.A(\reg_temp[155] ),
    .B(net549),
    .X(net324));
 sky130_fd_sc_hd__and2_1 _1798_ (.A(\reg_temp[156] ),
    .B(net549),
    .X(net325));
 sky130_fd_sc_hd__and2_1 _1799_ (.A(\reg_temp[157] ),
    .B(net550),
    .X(net326));
 sky130_fd_sc_hd__and2_1 _1800_ (.A(\reg_temp[158] ),
    .B(net550),
    .X(net327));
 sky130_fd_sc_hd__and2_1 _1801_ (.A(\reg_temp[159] ),
    .B(net550),
    .X(net328));
 sky130_fd_sc_hd__and2_1 _1802_ (.A(\reg_temp[160] ),
    .B(net550),
    .X(net330));
 sky130_fd_sc_hd__and2_1 _1803_ (.A(\reg_temp[161] ),
    .B(net545),
    .X(net331));
 sky130_fd_sc_hd__and2_1 _1804_ (.A(\reg_temp[162] ),
    .B(net545),
    .X(net332));
 sky130_fd_sc_hd__or3b_1 _1805_ (.A(_0570_),
    .B(net179),
    .C_N(net178),
    .X(_0947_));
 sky130_fd_sc_hd__or4b_1 _1806_ (.A(net177),
    .B(net189),
    .C(_0947_),
    .D_N(net176),
    .X(_0948_));
 sky130_fd_sc_hd__nor2_1 _1807_ (.A(_0942_),
    .B(_0948_),
    .Y(_0003_));
 sky130_fd_sc_hd__or4_1 _1808_ (.A(net174),
    .B(net173),
    .C(net176),
    .D(net177),
    .X(_0949_));
 sky130_fd_sc_hd__or3b_1 _1809_ (.A(_0949_),
    .B(net179),
    .C_N(net178),
    .X(_0950_));
 sky130_fd_sc_hd__or4_1 _1810_ (.A(net172),
    .B(_0521_),
    .C(_0524_),
    .D(_0950_),
    .X(_0951_));
 sky130_fd_sc_hd__nor2_1 _1811_ (.A(_0573_),
    .B(_0951_),
    .Y(_0000_));
 sky130_fd_sc_hd__and3_1 _1812_ (.A(\reg_temp[0] ),
    .B(\current_state[0] ),
    .C(\current_state[1] ),
    .X(net426));
 sky130_fd_sc_hd__clkbuf_1 _1813_ (.A(\current_state[1] ),
    .X(_0005_));
 sky130_fd_sc_hd__inv_2 _1814_ (.A(net598),
    .Y(_0009_));
 sky130_fd_sc_hd__inv_2 _1815_ (.A(net598),
    .Y(_0010_));
 sky130_fd_sc_hd__inv_2 _1816_ (.A(net598),
    .Y(_0011_));
 sky130_fd_sc_hd__inv_2 _1817_ (.A(net600),
    .Y(_0012_));
 sky130_fd_sc_hd__inv_2 _1818_ (.A(net600),
    .Y(_0013_));
 sky130_fd_sc_hd__inv_2 _1819_ (.A(net600),
    .Y(_0014_));
 sky130_fd_sc_hd__inv_2 _1820_ (.A(net600),
    .Y(_0015_));
 sky130_fd_sc_hd__inv_2 _1821_ (.A(net600),
    .Y(_0016_));
 sky130_fd_sc_hd__inv_2 _1822_ (.A(net598),
    .Y(_0017_));
 sky130_fd_sc_hd__inv_2 _1823_ (.A(net598),
    .Y(_0018_));
 sky130_fd_sc_hd__inv_2 _1824_ (.A(net598),
    .Y(_0019_));
 sky130_fd_sc_hd__inv_2 _1825_ (.A(net600),
    .Y(_0020_));
 sky130_fd_sc_hd__inv_2 _1826_ (.A(net600),
    .Y(_0021_));
 sky130_fd_sc_hd__inv_2 _1827_ (.A(net600),
    .Y(_0022_));
 sky130_fd_sc_hd__inv_2 _1828_ (.A(net600),
    .Y(_0023_));
 sky130_fd_sc_hd__inv_2 _1829_ (.A(net600),
    .Y(_0024_));
 sky130_fd_sc_hd__inv_2 _1830_ (.A(net600),
    .Y(_0025_));
 sky130_fd_sc_hd__inv_2 _1831_ (.A(net600),
    .Y(_0026_));
 sky130_fd_sc_hd__inv_2 _1832_ (.A(net602),
    .Y(_0027_));
 sky130_fd_sc_hd__inv_2 _1833_ (.A(net602),
    .Y(_0028_));
 sky130_fd_sc_hd__inv_2 _1834_ (.A(net602),
    .Y(_0029_));
 sky130_fd_sc_hd__inv_2 _1835_ (.A(net602),
    .Y(_0030_));
 sky130_fd_sc_hd__inv_2 _1836_ (.A(net600),
    .Y(_0031_));
 sky130_fd_sc_hd__inv_2 _1837_ (.A(net600),
    .Y(_0032_));
 sky130_fd_sc_hd__inv_2 _1838_ (.A(net600),
    .Y(_0033_));
 sky130_fd_sc_hd__inv_2 _1839_ (.A(net602),
    .Y(_0034_));
 sky130_fd_sc_hd__inv_2 _1840_ (.A(net602),
    .Y(_0035_));
 sky130_fd_sc_hd__inv_2 _1841_ (.A(net602),
    .Y(_0036_));
 sky130_fd_sc_hd__inv_2 _1842_ (.A(net601),
    .Y(_0037_));
 sky130_fd_sc_hd__inv_2 _1843_ (.A(net601),
    .Y(_0038_));
 sky130_fd_sc_hd__inv_2 _1844_ (.A(net601),
    .Y(_0039_));
 sky130_fd_sc_hd__inv_2 _1845_ (.A(net601),
    .Y(_0040_));
 sky130_fd_sc_hd__inv_2 _1846_ (.A(net601),
    .Y(_0041_));
 sky130_fd_sc_hd__inv_2 _1847_ (.A(net601),
    .Y(_0042_));
 sky130_fd_sc_hd__inv_2 _1848_ (.A(net601),
    .Y(_0043_));
 sky130_fd_sc_hd__inv_2 _1849_ (.A(net601),
    .Y(_0044_));
 sky130_fd_sc_hd__inv_2 _1850_ (.A(net601),
    .Y(_0045_));
 sky130_fd_sc_hd__inv_2 _1851_ (.A(net601),
    .Y(_0046_));
 sky130_fd_sc_hd__inv_2 _1852_ (.A(net600),
    .Y(_0047_));
 sky130_fd_sc_hd__inv_2 _1853_ (.A(net598),
    .Y(_0048_));
 sky130_fd_sc_hd__inv_2 _1854_ (.A(net598),
    .Y(_0049_));
 sky130_fd_sc_hd__inv_2 _1855_ (.A(net598),
    .Y(_0050_));
 sky130_fd_sc_hd__inv_2 _1856_ (.A(net599),
    .Y(_0051_));
 sky130_fd_sc_hd__inv_2 _1857_ (.A(net599),
    .Y(_0052_));
 sky130_fd_sc_hd__inv_2 _1858_ (.A(net606),
    .Y(_0053_));
 sky130_fd_sc_hd__inv_2 _1859_ (.A(net606),
    .Y(_0054_));
 sky130_fd_sc_hd__inv_2 _1860_ (.A(net606),
    .Y(_0055_));
 sky130_fd_sc_hd__inv_2 _1861_ (.A(net603),
    .Y(_0056_));
 sky130_fd_sc_hd__inv_2 _1862_ (.A(net603),
    .Y(_0057_));
 sky130_fd_sc_hd__inv_2 _1863_ (.A(net603),
    .Y(_0058_));
 sky130_fd_sc_hd__inv_2 _1864_ (.A(net604),
    .Y(_0059_));
 sky130_fd_sc_hd__inv_2 _1865_ (.A(net604),
    .Y(_0060_));
 sky130_fd_sc_hd__inv_2 _1866_ (.A(net604),
    .Y(_0061_));
 sky130_fd_sc_hd__inv_2 _1867_ (.A(net604),
    .Y(_0062_));
 sky130_fd_sc_hd__inv_2 _1868_ (.A(net604),
    .Y(_0063_));
 sky130_fd_sc_hd__inv_2 _1869_ (.A(net610),
    .Y(_0064_));
 sky130_fd_sc_hd__inv_2 _1870_ (.A(net610),
    .Y(_0065_));
 sky130_fd_sc_hd__inv_2 _1871_ (.A(net610),
    .Y(_0066_));
 sky130_fd_sc_hd__inv_2 _1872_ (.A(net610),
    .Y(_0067_));
 sky130_fd_sc_hd__inv_2 _1873_ (.A(net610),
    .Y(_0068_));
 sky130_fd_sc_hd__inv_2 _1874_ (.A(net610),
    .Y(_0069_));
 sky130_fd_sc_hd__inv_2 _1875_ (.A(net610),
    .Y(_0070_));
 sky130_fd_sc_hd__inv_2 _1876_ (.A(net610),
    .Y(_0071_));
 sky130_fd_sc_hd__inv_2 _1877_ (.A(net617),
    .Y(_0072_));
 sky130_fd_sc_hd__inv_2 _1878_ (.A(net617),
    .Y(_0073_));
 sky130_fd_sc_hd__inv_2 _1879_ (.A(net612),
    .Y(_0074_));
 sky130_fd_sc_hd__inv_2 _1880_ (.A(net613),
    .Y(_0075_));
 sky130_fd_sc_hd__inv_2 _1881_ (.A(net616),
    .Y(_0076_));
 sky130_fd_sc_hd__inv_2 _1882_ (.A(net616),
    .Y(_0077_));
 sky130_fd_sc_hd__inv_2 _1883_ (.A(net616),
    .Y(_0078_));
 sky130_fd_sc_hd__inv_2 _1884_ (.A(net617),
    .Y(_0079_));
 sky130_fd_sc_hd__inv_2 _1885_ (.A(net617),
    .Y(_0080_));
 sky130_fd_sc_hd__inv_2 _1886_ (.A(net616),
    .Y(_0081_));
 sky130_fd_sc_hd__inv_2 _1887_ (.A(net616),
    .Y(_0082_));
 sky130_fd_sc_hd__inv_2 _1888_ (.A(net617),
    .Y(_0083_));
 sky130_fd_sc_hd__inv_2 _1889_ (.A(net617),
    .Y(_0084_));
 sky130_fd_sc_hd__inv_2 _1890_ (.A(net616),
    .Y(_0085_));
 sky130_fd_sc_hd__inv_2 _1891_ (.A(net614),
    .Y(_0086_));
 sky130_fd_sc_hd__inv_2 _1892_ (.A(net614),
    .Y(_0087_));
 sky130_fd_sc_hd__inv_2 _1893_ (.A(net614),
    .Y(_0088_));
 sky130_fd_sc_hd__inv_2 _1894_ (.A(net606),
    .Y(_0089_));
 sky130_fd_sc_hd__inv_2 _1895_ (.A(net613),
    .Y(_0090_));
 sky130_fd_sc_hd__inv_2 _1896_ (.A(net613),
    .Y(_0091_));
 sky130_fd_sc_hd__inv_2 _1897_ (.A(net612),
    .Y(_0092_));
 sky130_fd_sc_hd__inv_2 _1898_ (.A(net606),
    .Y(_0093_));
 sky130_fd_sc_hd__inv_2 _1899_ (.A(net606),
    .Y(_0094_));
 sky130_fd_sc_hd__inv_2 _1900_ (.A(net599),
    .Y(_0095_));
 sky130_fd_sc_hd__inv_2 _1901_ (.A(net606),
    .Y(_0096_));
 sky130_fd_sc_hd__inv_2 _1902_ (.A(net599),
    .Y(_0097_));
 sky130_fd_sc_hd__inv_2 _1903_ (.A(net599),
    .Y(_0098_));
 sky130_fd_sc_hd__inv_2 _1904_ (.A(net599),
    .Y(_0099_));
 sky130_fd_sc_hd__inv_2 _1905_ (.A(net599),
    .Y(_0100_));
 sky130_fd_sc_hd__inv_2 _1906_ (.A(net601),
    .Y(_0101_));
 sky130_fd_sc_hd__inv_2 _1907_ (.A(net601),
    .Y(_0102_));
 sky130_fd_sc_hd__inv_2 _1908_ (.A(net602),
    .Y(_0103_));
 sky130_fd_sc_hd__inv_2 _1909_ (.A(net602),
    .Y(_0104_));
 sky130_fd_sc_hd__inv_2 _1910_ (.A(net601),
    .Y(_0105_));
 sky130_fd_sc_hd__inv_2 _1911_ (.A(net599),
    .Y(_0106_));
 sky130_fd_sc_hd__inv_2 _1912_ (.A(net599),
    .Y(_0107_));
 sky130_fd_sc_hd__inv_2 _1913_ (.A(net599),
    .Y(_0108_));
 sky130_fd_sc_hd__inv_2 _1914_ (.A(net601),
    .Y(_0109_));
 sky130_fd_sc_hd__inv_2 _1915_ (.A(net601),
    .Y(_0110_));
 sky130_fd_sc_hd__inv_2 _1916_ (.A(net601),
    .Y(_0111_));
 sky130_fd_sc_hd__inv_2 _1917_ (.A(net603),
    .Y(_0112_));
 sky130_fd_sc_hd__inv_2 _1918_ (.A(net603),
    .Y(_0113_));
 sky130_fd_sc_hd__inv_2 _1919_ (.A(net603),
    .Y(_0114_));
 sky130_fd_sc_hd__inv_2 _1920_ (.A(net602),
    .Y(_0115_));
 sky130_fd_sc_hd__inv_2 _1921_ (.A(net602),
    .Y(_0116_));
 sky130_fd_sc_hd__inv_2 _1922_ (.A(net602),
    .Y(_0117_));
 sky130_fd_sc_hd__inv_2 _1923_ (.A(net603),
    .Y(_0118_));
 sky130_fd_sc_hd__inv_2 _1924_ (.A(net603),
    .Y(_0119_));
 sky130_fd_sc_hd__inv_2 _1925_ (.A(net603),
    .Y(_0120_));
 sky130_fd_sc_hd__inv_2 _1926_ (.A(net603),
    .Y(_0121_));
 sky130_fd_sc_hd__inv_2 _1927_ (.A(net603),
    .Y(_0122_));
 sky130_fd_sc_hd__inv_2 _1928_ (.A(net603),
    .Y(_0123_));
 sky130_fd_sc_hd__inv_2 _1929_ (.A(net603),
    .Y(_0124_));
 sky130_fd_sc_hd__inv_2 _1930_ (.A(net603),
    .Y(_0125_));
 sky130_fd_sc_hd__inv_2 _1931_ (.A(net605),
    .Y(_0126_));
 sky130_fd_sc_hd__inv_2 _1932_ (.A(net604),
    .Y(_0127_));
 sky130_fd_sc_hd__inv_2 _1933_ (.A(net604),
    .Y(_0128_));
 sky130_fd_sc_hd__inv_2 _1934_ (.A(net604),
    .Y(_0129_));
 sky130_fd_sc_hd__inv_2 _1935_ (.A(net604),
    .Y(_0130_));
 sky130_fd_sc_hd__inv_2 _1936_ (.A(net605),
    .Y(_0131_));
 sky130_fd_sc_hd__inv_2 _1937_ (.A(net605),
    .Y(_0132_));
 sky130_fd_sc_hd__inv_2 _1938_ (.A(net604),
    .Y(_0133_));
 sky130_fd_sc_hd__inv_2 _1939_ (.A(net604),
    .Y(_0134_));
 sky130_fd_sc_hd__inv_2 _1940_ (.A(net603),
    .Y(_0135_));
 sky130_fd_sc_hd__inv_2 _1941_ (.A(net603),
    .Y(_0136_));
 sky130_fd_sc_hd__inv_2 _1942_ (.A(net606),
    .Y(_0137_));
 sky130_fd_sc_hd__inv_2 _1943_ (.A(net606),
    .Y(_0138_));
 sky130_fd_sc_hd__inv_2 _1944_ (.A(net606),
    .Y(_0139_));
 sky130_fd_sc_hd__inv_2 _1945_ (.A(net606),
    .Y(_0140_));
 sky130_fd_sc_hd__inv_2 _1946_ (.A(net606),
    .Y(_0141_));
 sky130_fd_sc_hd__inv_2 _1947_ (.A(net606),
    .Y(_0142_));
 sky130_fd_sc_hd__inv_2 _1948_ (.A(net606),
    .Y(_0143_));
 sky130_fd_sc_hd__inv_2 _1949_ (.A(net606),
    .Y(_0144_));
 sky130_fd_sc_hd__inv_2 _1950_ (.A(net604),
    .Y(_0145_));
 sky130_fd_sc_hd__inv_2 _1951_ (.A(net604),
    .Y(_0146_));
 sky130_fd_sc_hd__inv_2 _1952_ (.A(net604),
    .Y(_0147_));
 sky130_fd_sc_hd__inv_2 _1953_ (.A(net604),
    .Y(_0148_));
 sky130_fd_sc_hd__inv_2 _1954_ (.A(net604),
    .Y(_0149_));
 sky130_fd_sc_hd__inv_2 _1955_ (.A(net605),
    .Y(_0150_));
 sky130_fd_sc_hd__inv_2 _1956_ (.A(net605),
    .Y(_0151_));
 sky130_fd_sc_hd__inv_2 _1957_ (.A(net605),
    .Y(_0152_));
 sky130_fd_sc_hd__inv_2 _1958_ (.A(net610),
    .Y(_0153_));
 sky130_fd_sc_hd__inv_2 _1959_ (.A(net610),
    .Y(_0154_));
 sky130_fd_sc_hd__inv_2 _1960_ (.A(net610),
    .Y(_0155_));
 sky130_fd_sc_hd__inv_2 _1961_ (.A(net610),
    .Y(_0156_));
 sky130_fd_sc_hd__inv_2 _1962_ (.A(net610),
    .Y(_0157_));
 sky130_fd_sc_hd__inv_2 _1963_ (.A(net610),
    .Y(_0158_));
 sky130_fd_sc_hd__inv_2 _1964_ (.A(net611),
    .Y(_0159_));
 sky130_fd_sc_hd__inv_2 _1965_ (.A(net611),
    .Y(_0160_));
 sky130_fd_sc_hd__inv_2 _1966_ (.A(net617),
    .Y(_0161_));
 sky130_fd_sc_hd__inv_2 _1967_ (.A(net616),
    .Y(_0162_));
 sky130_fd_sc_hd__inv_2 _1968_ (.A(net614),
    .Y(_0163_));
 sky130_fd_sc_hd__inv_2 _1969_ (.A(net614),
    .Y(_0164_));
 sky130_fd_sc_hd__inv_2 _1970_ (.A(net616),
    .Y(_0165_));
 sky130_fd_sc_hd__inv_2 _1971_ (.A(net616),
    .Y(_0166_));
 sky130_fd_sc_hd__inv_2 _1972_ (.A(net616),
    .Y(_0167_));
 sky130_fd_sc_hd__inv_2 _1973_ (.A(net616),
    .Y(_0168_));
 sky130_fd_sc_hd__inv_2 _1974_ (.A(net616),
    .Y(_0169_));
 sky130_fd_sc_hd__inv_2 _1975_ (.A(net616),
    .Y(_0170_));
 sky130_fd_sc_hd__inv_2 _1976_ (.A(net616),
    .Y(_0171_));
 sky130_fd_sc_hd__inv_2 _1977_ (.A(net616),
    .Y(_0172_));
 sky130_fd_sc_hd__inv_2 _1978_ (.A(net617),
    .Y(_0173_));
 sky130_fd_sc_hd__inv_2 _1979_ (.A(net616),
    .Y(_0174_));
 sky130_fd_sc_hd__inv_2 _1980_ (.A(net614),
    .Y(_0175_));
 sky130_fd_sc_hd__inv_2 _1981_ (.A(net614),
    .Y(_0176_));
 sky130_fd_sc_hd__inv_2 _1982_ (.A(net614),
    .Y(_0177_));
 sky130_fd_sc_hd__inv_2 _1983_ (.A(net598),
    .Y(_0178_));
 sky130_fd_sc_hd__inv_2 _1984_ (.A(net598),
    .Y(_0179_));
 sky130_fd_sc_hd__inv_2 _1985_ (.A(net598),
    .Y(_0180_));
 sky130_fd_sc_hd__inv_2 _1986_ (.A(net598),
    .Y(_0181_));
 sky130_fd_sc_hd__inv_2 _1987_ (.A(net598),
    .Y(_0182_));
 sky130_fd_sc_hd__inv_2 _1988_ (.A(net598),
    .Y(_0183_));
 sky130_fd_sc_hd__inv_2 _1989_ (.A(net607),
    .Y(_0184_));
 sky130_fd_sc_hd__inv_2 _1990_ (.A(net607),
    .Y(_0185_));
 sky130_fd_sc_hd__inv_2 _1991_ (.A(net607),
    .Y(_0186_));
 sky130_fd_sc_hd__inv_2 _1992_ (.A(net607),
    .Y(_0187_));
 sky130_fd_sc_hd__inv_2 _1993_ (.A(net607),
    .Y(_0188_));
 sky130_fd_sc_hd__inv_2 _1994_ (.A(net607),
    .Y(_0189_));
 sky130_fd_sc_hd__inv_2 _1995_ (.A(net610),
    .Y(_0190_));
 sky130_fd_sc_hd__inv_2 _1996_ (.A(net607),
    .Y(_0191_));
 sky130_fd_sc_hd__inv_2 _1997_ (.A(net607),
    .Y(_0192_));
 sky130_fd_sc_hd__inv_2 _1998_ (.A(net607),
    .Y(_0193_));
 sky130_fd_sc_hd__inv_2 _1999_ (.A(net607),
    .Y(_0194_));
 sky130_fd_sc_hd__inv_2 _2000_ (.A(net607),
    .Y(_0195_));
 sky130_fd_sc_hd__inv_2 _2001_ (.A(net607),
    .Y(_0196_));
 sky130_fd_sc_hd__inv_2 _2002_ (.A(net610),
    .Y(_0197_));
 sky130_fd_sc_hd__inv_2 _2003_ (.A(net607),
    .Y(_0198_));
 sky130_fd_sc_hd__inv_2 _2004_ (.A(net607),
    .Y(_0199_));
 sky130_fd_sc_hd__inv_2 _2005_ (.A(net609),
    .Y(_0200_));
 sky130_fd_sc_hd__inv_2 _2006_ (.A(net607),
    .Y(_0201_));
 sky130_fd_sc_hd__inv_2 _2007_ (.A(net611),
    .Y(_0202_));
 sky130_fd_sc_hd__inv_2 _2008_ (.A(net607),
    .Y(_0203_));
 sky130_fd_sc_hd__inv_2 _2009_ (.A(net609),
    .Y(_0204_));
 sky130_fd_sc_hd__inv_2 _2010_ (.A(net608),
    .Y(_0205_));
 sky130_fd_sc_hd__inv_2 _2011_ (.A(net609),
    .Y(_0206_));
 sky130_fd_sc_hd__inv_2 _2012_ (.A(net608),
    .Y(_0207_));
 sky130_fd_sc_hd__inv_2 _2013_ (.A(net608),
    .Y(_0208_));
 sky130_fd_sc_hd__inv_2 _2014_ (.A(net608),
    .Y(_0209_));
 sky130_fd_sc_hd__inv_2 _2015_ (.A(net608),
    .Y(_0210_));
 sky130_fd_sc_hd__inv_2 _2016_ (.A(net609),
    .Y(_0211_));
 sky130_fd_sc_hd__inv_2 _2017_ (.A(net611),
    .Y(_0212_));
 sky130_fd_sc_hd__inv_2 _2018_ (.A(net608),
    .Y(_0213_));
 sky130_fd_sc_hd__inv_2 _2019_ (.A(net608),
    .Y(_0214_));
 sky130_fd_sc_hd__inv_2 _2020_ (.A(net608),
    .Y(_0215_));
 sky130_fd_sc_hd__inv_2 _2021_ (.A(net609),
    .Y(_0216_));
 sky130_fd_sc_hd__inv_2 _2022_ (.A(net611),
    .Y(_0217_));
 sky130_fd_sc_hd__inv_2 _2023_ (.A(net608),
    .Y(_0218_));
 sky130_fd_sc_hd__inv_2 _2024_ (.A(net608),
    .Y(_0219_));
 sky130_fd_sc_hd__inv_2 _2025_ (.A(net611),
    .Y(_0220_));
 sky130_fd_sc_hd__inv_2 _2026_ (.A(net611),
    .Y(_0221_));
 sky130_fd_sc_hd__inv_2 _2027_ (.A(net609),
    .Y(_0222_));
 sky130_fd_sc_hd__inv_2 _2028_ (.A(net608),
    .Y(_0223_));
 sky130_fd_sc_hd__inv_2 _2029_ (.A(net608),
    .Y(_0224_));
 sky130_fd_sc_hd__inv_2 _2030_ (.A(net608),
    .Y(_0225_));
 sky130_fd_sc_hd__inv_2 _2031_ (.A(net608),
    .Y(_0226_));
 sky130_fd_sc_hd__inv_2 _2032_ (.A(net608),
    .Y(_0227_));
 sky130_fd_sc_hd__inv_2 _2033_ (.A(net608),
    .Y(_0228_));
 sky130_fd_sc_hd__inv_2 _2034_ (.A(net609),
    .Y(_0229_));
 sky130_fd_sc_hd__inv_2 _2035_ (.A(net612),
    .Y(_0230_));
 sky130_fd_sc_hd__inv_2 _2036_ (.A(net612),
    .Y(_0231_));
 sky130_fd_sc_hd__inv_2 _2037_ (.A(net612),
    .Y(_0232_));
 sky130_fd_sc_hd__inv_2 _2038_ (.A(net615),
    .Y(_0233_));
 sky130_fd_sc_hd__inv_2 _2039_ (.A(net617),
    .Y(_0234_));
 sky130_fd_sc_hd__inv_2 _2040_ (.A(net612),
    .Y(_0235_));
 sky130_fd_sc_hd__inv_2 _2041_ (.A(net615),
    .Y(_0236_));
 sky130_fd_sc_hd__inv_2 _2042_ (.A(net612),
    .Y(_0237_));
 sky130_fd_sc_hd__inv_2 _2043_ (.A(net612),
    .Y(_0238_));
 sky130_fd_sc_hd__inv_2 _2044_ (.A(net612),
    .Y(_0239_));
 sky130_fd_sc_hd__inv_2 _2045_ (.A(net612),
    .Y(_0240_));
 sky130_fd_sc_hd__inv_2 _2046_ (.A(net612),
    .Y(_0241_));
 sky130_fd_sc_hd__inv_2 _2047_ (.A(net612),
    .Y(_0242_));
 sky130_fd_sc_hd__inv_2 _2048_ (.A(net615),
    .Y(_0243_));
 sky130_fd_sc_hd__inv_2 _2049_ (.A(net615),
    .Y(_0244_));
 sky130_fd_sc_hd__inv_2 _2050_ (.A(net612),
    .Y(_0245_));
 sky130_fd_sc_hd__inv_2 _2051_ (.A(net612),
    .Y(_0246_));
 sky130_fd_sc_hd__inv_2 _2052_ (.A(net615),
    .Y(_0247_));
 sky130_fd_sc_hd__inv_2 _2053_ (.A(net612),
    .Y(_0248_));
 sky130_fd_sc_hd__inv_2 _2054_ (.A(net615),
    .Y(_0249_));
 sky130_fd_sc_hd__inv_2 _2055_ (.A(net613),
    .Y(_0250_));
 sky130_fd_sc_hd__inv_2 _2056_ (.A(net613),
    .Y(_0251_));
 sky130_fd_sc_hd__inv_2 _2057_ (.A(net613),
    .Y(_0252_));
 sky130_fd_sc_hd__inv_2 _2058_ (.A(net613),
    .Y(_0253_));
 sky130_fd_sc_hd__inv_2 _2059_ (.A(net613),
    .Y(_0254_));
 sky130_fd_sc_hd__inv_2 _2060_ (.A(net613),
    .Y(_0255_));
 sky130_fd_sc_hd__inv_2 _2061_ (.A(net615),
    .Y(_0256_));
 sky130_fd_sc_hd__inv_2 _2062_ (.A(net613),
    .Y(_0257_));
 sky130_fd_sc_hd__inv_2 _2063_ (.A(net613),
    .Y(_0258_));
 sky130_fd_sc_hd__inv_2 _2064_ (.A(net613),
    .Y(_0259_));
 sky130_fd_sc_hd__inv_2 _2065_ (.A(net612),
    .Y(_0260_));
 sky130_fd_sc_hd__inv_2 _2066_ (.A(net613),
    .Y(_0261_));
 sky130_fd_sc_hd__inv_2 _2067_ (.A(net613),
    .Y(_0262_));
 sky130_fd_sc_hd__inv_2 _2068_ (.A(net613),
    .Y(_0263_));
 sky130_fd_sc_hd__inv_2 _2069_ (.A(net613),
    .Y(_0264_));
 sky130_fd_sc_hd__dfrtp_4 _2070_ (.CLK(clknet_leaf_26_wb_clk_i),
    .D(net708),
    .RESET_B(_0008_),
    .Q(\reg_temp[0] ));
 sky130_fd_sc_hd__dfrtp_4 _2071_ (.CLK(clknet_leaf_26_wb_clk_i),
    .D(net690),
    .RESET_B(_0009_),
    .Q(\reg_temp[1] ));
 sky130_fd_sc_hd__dfrtp_4 _2072_ (.CLK(clknet_leaf_26_wb_clk_i),
    .D(net676),
    .RESET_B(_0010_),
    .Q(\reg_temp[2] ));
 sky130_fd_sc_hd__dfrtp_4 _2073_ (.CLK(clknet_leaf_26_wb_clk_i),
    .D(_0268_),
    .RESET_B(_0011_),
    .Q(\reg_temp[3] ));
 sky130_fd_sc_hd__dfrtp_4 _2074_ (.CLK(clknet_leaf_3_wb_clk_i),
    .D(net1609),
    .RESET_B(_0012_),
    .Q(\reg_temp[4] ));
 sky130_fd_sc_hd__dfrtp_4 _2075_ (.CLK(clknet_leaf_3_wb_clk_i),
    .D(_0270_),
    .RESET_B(_0013_),
    .Q(\reg_temp[5] ));
 sky130_fd_sc_hd__dfrtp_4 _2076_ (.CLK(clknet_leaf_4_wb_clk_i),
    .D(net739),
    .RESET_B(_0014_),
    .Q(\reg_temp[6] ));
 sky130_fd_sc_hd__dfrtp_4 _2077_ (.CLK(clknet_leaf_5_wb_clk_i),
    .D(net1575),
    .RESET_B(_0015_),
    .Q(\reg_temp[7] ));
 sky130_fd_sc_hd__dfrtp_4 _2078_ (.CLK(clknet_leaf_3_wb_clk_i),
    .D(_0273_),
    .RESET_B(_0016_),
    .Q(\reg_temp[8] ));
 sky130_fd_sc_hd__dfrtp_4 _2079_ (.CLK(clknet_leaf_26_wb_clk_i),
    .D(net760),
    .RESET_B(_0017_),
    .Q(\reg_temp[9] ));
 sky130_fd_sc_hd__dfrtp_4 _2080_ (.CLK(clknet_leaf_26_wb_clk_i),
    .D(net713),
    .RESET_B(_0018_),
    .Q(\reg_temp[10] ));
 sky130_fd_sc_hd__dfrtp_4 _2081_ (.CLK(clknet_leaf_26_wb_clk_i),
    .D(net815),
    .RESET_B(_0019_),
    .Q(\reg_temp[11] ));
 sky130_fd_sc_hd__dfrtp_4 _2082_ (.CLK(clknet_leaf_3_wb_clk_i),
    .D(_0277_),
    .RESET_B(_0020_),
    .Q(\reg_temp[12] ));
 sky130_fd_sc_hd__dfrtp_4 _2083_ (.CLK(clknet_leaf_3_wb_clk_i),
    .D(_0278_),
    .RESET_B(_0021_),
    .Q(\reg_temp[13] ));
 sky130_fd_sc_hd__dfrtp_4 _2084_ (.CLK(clknet_leaf_3_wb_clk_i),
    .D(net1547),
    .RESET_B(_0022_),
    .Q(\reg_temp[14] ));
 sky130_fd_sc_hd__dfrtp_4 _2085_ (.CLK(clknet_leaf_3_wb_clk_i),
    .D(net1600),
    .RESET_B(_0023_),
    .Q(\reg_temp[15] ));
 sky130_fd_sc_hd__dfrtp_4 _2086_ (.CLK(clknet_leaf_4_wb_clk_i),
    .D(net1431),
    .RESET_B(_0024_),
    .Q(\reg_temp[16] ));
 sky130_fd_sc_hd__dfrtp_4 _2087_ (.CLK(clknet_leaf_4_wb_clk_i),
    .D(_0282_),
    .RESET_B(_0025_),
    .Q(\reg_temp[17] ));
 sky130_fd_sc_hd__dfrtp_4 _2088_ (.CLK(clknet_leaf_4_wb_clk_i),
    .D(_0283_),
    .RESET_B(_0026_),
    .Q(\reg_temp[18] ));
 sky130_fd_sc_hd__dfrtp_4 _2089_ (.CLK(clknet_leaf_5_wb_clk_i),
    .D(_0284_),
    .RESET_B(_0027_),
    .Q(\reg_temp[19] ));
 sky130_fd_sc_hd__dfrtp_4 _2090_ (.CLK(clknet_leaf_5_wb_clk_i),
    .D(_0285_),
    .RESET_B(_0028_),
    .Q(\reg_temp[20] ));
 sky130_fd_sc_hd__dfrtp_4 _2091_ (.CLK(clknet_leaf_5_wb_clk_i),
    .D(_0286_),
    .RESET_B(_0029_),
    .Q(\reg_temp[21] ));
 sky130_fd_sc_hd__dfrtp_4 _2092_ (.CLK(clknet_leaf_5_wb_clk_i),
    .D(_0287_),
    .RESET_B(_0030_),
    .Q(\reg_temp[22] ));
 sky130_fd_sc_hd__dfrtp_4 _2093_ (.CLK(clknet_leaf_3_wb_clk_i),
    .D(_0288_),
    .RESET_B(_0031_),
    .Q(\reg_temp[23] ));
 sky130_fd_sc_hd__dfrtp_4 _2094_ (.CLK(clknet_leaf_3_wb_clk_i),
    .D(net1585),
    .RESET_B(_0032_),
    .Q(\reg_temp[24] ));
 sky130_fd_sc_hd__dfrtp_4 _2095_ (.CLK(clknet_leaf_3_wb_clk_i),
    .D(_0290_),
    .RESET_B(_0033_),
    .Q(\reg_temp[25] ));
 sky130_fd_sc_hd__dfrtp_4 _2096_ (.CLK(clknet_leaf_4_wb_clk_i),
    .D(net1596),
    .RESET_B(_0034_),
    .Q(\reg_temp[26] ));
 sky130_fd_sc_hd__dfrtp_4 _2097_ (.CLK(clknet_leaf_4_wb_clk_i),
    .D(_0292_),
    .RESET_B(_0035_),
    .Q(\reg_temp[27] ));
 sky130_fd_sc_hd__dfrtp_4 _2098_ (.CLK(clknet_leaf_4_wb_clk_i),
    .D(_0293_),
    .RESET_B(_0036_),
    .Q(\reg_temp[28] ));
 sky130_fd_sc_hd__dfrtp_4 _2099_ (.CLK(clknet_leaf_5_wb_clk_i),
    .D(_0294_),
    .RESET_B(_0037_),
    .Q(\reg_temp[29] ));
 sky130_fd_sc_hd__dfrtp_4 _2100_ (.CLK(clknet_leaf_5_wb_clk_i),
    .D(_0295_),
    .RESET_B(_0038_),
    .Q(\reg_temp[30] ));
 sky130_fd_sc_hd__dfrtp_4 _2101_ (.CLK(clknet_leaf_5_wb_clk_i),
    .D(_0296_),
    .RESET_B(_0039_),
    .Q(\reg_temp[31] ));
 sky130_fd_sc_hd__dfrtp_4 _2102_ (.CLK(clknet_leaf_5_wb_clk_i),
    .D(_0297_),
    .RESET_B(_0040_),
    .Q(\reg_temp[32] ));
 sky130_fd_sc_hd__dfrtp_4 _2103_ (.CLK(clknet_leaf_6_wb_clk_i),
    .D(net1591),
    .RESET_B(_0041_),
    .Q(\reg_temp[33] ));
 sky130_fd_sc_hd__dfrtp_4 _2104_ (.CLK(clknet_leaf_4_wb_clk_i),
    .D(_0299_),
    .RESET_B(_0042_),
    .Q(\reg_temp[34] ));
 sky130_fd_sc_hd__dfrtp_4 _2105_ (.CLK(clknet_leaf_4_wb_clk_i),
    .D(_0300_),
    .RESET_B(_0043_),
    .Q(\reg_temp[35] ));
 sky130_fd_sc_hd__dfrtp_4 _2106_ (.CLK(clknet_leaf_3_wb_clk_i),
    .D(_0301_),
    .RESET_B(_0044_),
    .Q(\reg_temp[36] ));
 sky130_fd_sc_hd__dfrtp_4 _2107_ (.CLK(clknet_leaf_2_wb_clk_i),
    .D(net1545),
    .RESET_B(_0045_),
    .Q(\reg_temp[37] ));
 sky130_fd_sc_hd__dfrtp_4 _2108_ (.CLK(clknet_leaf_2_wb_clk_i),
    .D(_0303_),
    .RESET_B(_0046_),
    .Q(\reg_temp[38] ));
 sky130_fd_sc_hd__dfrtp_4 _2109_ (.CLK(clknet_leaf_2_wb_clk_i),
    .D(_0304_),
    .RESET_B(_0047_),
    .Q(\reg_temp[39] ));
 sky130_fd_sc_hd__dfrtp_4 _2110_ (.CLK(clknet_leaf_26_wb_clk_i),
    .D(_0305_),
    .RESET_B(_0048_),
    .Q(\reg_temp[40] ));
 sky130_fd_sc_hd__dfrtp_4 _2111_ (.CLK(clknet_leaf_26_wb_clk_i),
    .D(_0306_),
    .RESET_B(_0049_),
    .Q(\reg_temp[41] ));
 sky130_fd_sc_hd__dfrtp_4 _2112_ (.CLK(clknet_leaf_26_wb_clk_i),
    .D(net1539),
    .RESET_B(_0050_),
    .Q(\reg_temp[42] ));
 sky130_fd_sc_hd__dfrtp_4 _2113_ (.CLK(clknet_leaf_26_wb_clk_i),
    .D(_0308_),
    .RESET_B(_0051_),
    .Q(\reg_temp[43] ));
 sky130_fd_sc_hd__dfrtp_4 _2114_ (.CLK(clknet_leaf_0_wb_clk_i),
    .D(net1515),
    .RESET_B(_0052_),
    .Q(\reg_temp[44] ));
 sky130_fd_sc_hd__dfrtp_4 _2115_ (.CLK(clknet_leaf_0_wb_clk_i),
    .D(net771),
    .RESET_B(_0053_),
    .Q(\reg_temp[45] ));
 sky130_fd_sc_hd__dfrtp_4 _2116_ (.CLK(clknet_leaf_0_wb_clk_i),
    .D(net857),
    .RESET_B(_0054_),
    .Q(\reg_temp[46] ));
 sky130_fd_sc_hd__dfrtp_4 _2117_ (.CLK(clknet_leaf_0_wb_clk_i),
    .D(net818),
    .RESET_B(_0055_),
    .Q(\reg_temp[47] ));
 sky130_fd_sc_hd__dfrtp_4 _2118_ (.CLK(clknet_leaf_1_wb_clk_i),
    .D(net809),
    .RESET_B(_0056_),
    .Q(\reg_temp[48] ));
 sky130_fd_sc_hd__dfrtp_4 _2119_ (.CLK(clknet_leaf_1_wb_clk_i),
    .D(_0314_),
    .RESET_B(_0057_),
    .Q(\reg_temp[49] ));
 sky130_fd_sc_hd__dfrtp_4 _2120_ (.CLK(clknet_leaf_1_wb_clk_i),
    .D(net836),
    .RESET_B(_0058_),
    .Q(\reg_temp[50] ));
 sky130_fd_sc_hd__dfrtp_4 _2121_ (.CLK(clknet_leaf_9_wb_clk_i),
    .D(net977),
    .RESET_B(_0059_),
    .Q(\reg_temp[51] ));
 sky130_fd_sc_hd__dfrtp_2 _2122_ (.CLK(clknet_leaf_8_wb_clk_i),
    .D(net950),
    .RESET_B(_0060_),
    .Q(\reg_temp[52] ));
 sky130_fd_sc_hd__dfrtp_2 _2123_ (.CLK(clknet_leaf_7_wb_clk_i),
    .D(net1023),
    .RESET_B(_0061_),
    .Q(\reg_temp[53] ));
 sky130_fd_sc_hd__dfrtp_2 _2124_ (.CLK(clknet_leaf_7_wb_clk_i),
    .D(net1060),
    .RESET_B(_0062_),
    .Q(\reg_temp[54] ));
 sky130_fd_sc_hd__dfrtp_2 _2125_ (.CLK(clknet_leaf_7_wb_clk_i),
    .D(net1050),
    .RESET_B(_0063_),
    .Q(\reg_temp[55] ));
 sky130_fd_sc_hd__dfrtp_4 _2126_ (.CLK(clknet_leaf_11_wb_clk_i),
    .D(net1110),
    .RESET_B(_0064_),
    .Q(\reg_temp[56] ));
 sky130_fd_sc_hd__dfrtp_4 _2127_ (.CLK(clknet_leaf_8_wb_clk_i),
    .D(net1603),
    .RESET_B(_0065_),
    .Q(\reg_temp[57] ));
 sky130_fd_sc_hd__dfrtp_2 _2128_ (.CLK(clknet_leaf_9_wb_clk_i),
    .D(net1129),
    .RESET_B(_0066_),
    .Q(\reg_temp[58] ));
 sky130_fd_sc_hd__dfrtp_2 _2129_ (.CLK(clknet_leaf_10_wb_clk_i),
    .D(net1122),
    .RESET_B(_0067_),
    .Q(\reg_temp[59] ));
 sky130_fd_sc_hd__dfrtp_2 _2130_ (.CLK(clknet_leaf_11_wb_clk_i),
    .D(net1163),
    .RESET_B(_0068_),
    .Q(\reg_temp[60] ));
 sky130_fd_sc_hd__dfrtp_2 _2131_ (.CLK(clknet_leaf_11_wb_clk_i),
    .D(_0326_),
    .RESET_B(_0069_),
    .Q(\reg_temp[61] ));
 sky130_fd_sc_hd__dfrtp_1 _2132_ (.CLK(clknet_leaf_12_wb_clk_i),
    .D(net966),
    .RESET_B(_0070_),
    .Q(\reg_temp[62] ));
 sky130_fd_sc_hd__dfrtp_1 _2133_ (.CLK(clknet_leaf_15_wb_clk_i),
    .D(net1134),
    .RESET_B(_0071_),
    .Q(\reg_temp[63] ));
 sky130_fd_sc_hd__dfrtp_1 _2134_ (.CLK(clknet_leaf_14_wb_clk_i),
    .D(net979),
    .RESET_B(_0072_),
    .Q(\reg_temp[64] ));
 sky130_fd_sc_hd__dfrtp_1 _2135_ (.CLK(clknet_leaf_14_wb_clk_i),
    .D(net990),
    .RESET_B(_0073_),
    .Q(\reg_temp[65] ));
 sky130_fd_sc_hd__dfrtp_1 _2136_ (.CLK(clknet_leaf_17_wb_clk_i),
    .D(net988),
    .RESET_B(_0074_),
    .Q(\reg_temp[66] ));
 sky130_fd_sc_hd__dfrtp_1 _2137_ (.CLK(clknet_leaf_18_wb_clk_i),
    .D(net1038),
    .RESET_B(_0075_),
    .Q(\reg_temp[67] ));
 sky130_fd_sc_hd__dfrtp_1 _2138_ (.CLK(clknet_leaf_14_wb_clk_i),
    .D(net1045),
    .RESET_B(_0076_),
    .Q(\reg_temp[68] ));
 sky130_fd_sc_hd__dfrtp_1 _2139_ (.CLK(clknet_leaf_14_wb_clk_i),
    .D(net1095),
    .RESET_B(_0077_),
    .Q(\reg_temp[69] ));
 sky130_fd_sc_hd__dfrtp_1 _2140_ (.CLK(clknet_leaf_14_wb_clk_i),
    .D(net1069),
    .RESET_B(_0078_),
    .Q(\reg_temp[70] ));
 sky130_fd_sc_hd__dfrtp_1 _2141_ (.CLK(clknet_leaf_13_wb_clk_i),
    .D(net1043),
    .RESET_B(_0079_),
    .Q(\reg_temp[71] ));
 sky130_fd_sc_hd__dfrtp_1 _2142_ (.CLK(clknet_leaf_12_wb_clk_i),
    .D(net1007),
    .RESET_B(_0080_),
    .Q(\reg_temp[72] ));
 sky130_fd_sc_hd__dfrtp_2 _2143_ (.CLK(clknet_leaf_13_wb_clk_i),
    .D(_0338_),
    .RESET_B(_0081_),
    .Q(\reg_temp[73] ));
 sky130_fd_sc_hd__dfrtp_1 _2144_ (.CLK(clknet_leaf_13_wb_clk_i),
    .D(net1117),
    .RESET_B(_0082_),
    .Q(\reg_temp[74] ));
 sky130_fd_sc_hd__dfrtp_2 _2145_ (.CLK(clknet_leaf_12_wb_clk_i),
    .D(_0340_),
    .RESET_B(_0083_),
    .Q(\reg_temp[75] ));
 sky130_fd_sc_hd__dfrtp_1 _2146_ (.CLK(clknet_leaf_12_wb_clk_i),
    .D(net1138),
    .RESET_B(_0084_),
    .Q(\reg_temp[76] ));
 sky130_fd_sc_hd__dfrtp_2 _2147_ (.CLK(clknet_leaf_14_wb_clk_i),
    .D(net957),
    .RESET_B(_0085_),
    .Q(\reg_temp[77] ));
 sky130_fd_sc_hd__dfrtp_1 _2148_ (.CLK(clknet_leaf_18_wb_clk_i),
    .D(net890),
    .RESET_B(_0086_),
    .Q(\reg_temp[78] ));
 sky130_fd_sc_hd__dfrtp_1 _2149_ (.CLK(clknet_leaf_18_wb_clk_i),
    .D(net828),
    .RESET_B(_0087_),
    .Q(\reg_temp[79] ));
 sky130_fd_sc_hd__dfrtp_1 _2150_ (.CLK(clknet_leaf_18_wb_clk_i),
    .D(net1082),
    .RESET_B(_0088_),
    .Q(\reg_temp[80] ));
 sky130_fd_sc_hd__dfrtp_4 _2151_ (.CLK(clknet_leaf_23_wb_clk_i),
    .D(net666),
    .RESET_B(_0089_),
    .Q(\reg_temp[81] ));
 sky130_fd_sc_hd__dfrtp_1 _2152_ (.CLK(clknet_leaf_20_wb_clk_i),
    .D(net1239),
    .RESET_B(_0090_),
    .Q(net445));
 sky130_fd_sc_hd__dfrtp_1 _2153_ (.CLK(clknet_leaf_20_wb_clk_i),
    .D(_0348_),
    .RESET_B(_0091_),
    .Q(net446));
 sky130_fd_sc_hd__dfrtp_1 _2154_ (.CLK(clknet_leaf_20_wb_clk_i),
    .D(net1090),
    .RESET_B(_0092_),
    .Q(net440));
 sky130_fd_sc_hd__dlxtn_1 _2155_ (.D(_0002_),
    .GATE_N(net591),
    .Q(net519));
 sky130_fd_sc_hd__dlxtn_1 _2156_ (.D(_0000_),
    .GATE_N(_0005_),
    .Q(enable_proc));
 sky130_fd_sc_hd__dfrtp_1 _2157_ (.CLK(clknet_leaf_24_wb_clk_i),
    .D(net781),
    .RESET_B(_0093_),
    .Q(net441));
 sky130_fd_sc_hd__dfrtp_1 _2158_ (.CLK(clknet_leaf_24_wb_clk_i),
    .D(net1146),
    .RESET_B(_0094_),
    .Q(net442));
 sky130_fd_sc_hd__dfrtp_1 _2159_ (.CLK(clknet_leaf_25_wb_clk_i),
    .D(net748),
    .RESET_B(_0095_),
    .Q(net443));
 sky130_fd_sc_hd__dfrtp_1 _2160_ (.CLK(clknet_leaf_24_wb_clk_i),
    .D(net1201),
    .RESET_B(_0096_),
    .Q(net444));
 sky130_fd_sc_hd__dlxtn_1 _2161_ (.D(_0001_),
    .GATE_N(_0006_),
    .Q(net515));
 sky130_fd_sc_hd__dfrtp_4 _2162_ (.CLK(clknet_leaf_0_wb_clk_i),
    .D(net1498),
    .RESET_B(_0097_),
    .Q(\reg_temp[82] ));
 sky130_fd_sc_hd__dfrtp_4 _2163_ (.CLK(clknet_leaf_26_wb_clk_i),
    .D(net698),
    .RESET_B(_0098_),
    .Q(\reg_temp[83] ));
 sky130_fd_sc_hd__dfrtp_4 _2164_ (.CLK(clknet_leaf_26_wb_clk_i),
    .D(net685),
    .RESET_B(_0099_),
    .Q(\reg_temp[84] ));
 sky130_fd_sc_hd__dfrtp_4 _2165_ (.CLK(clknet_leaf_0_wb_clk_i),
    .D(net1556),
    .RESET_B(_0100_),
    .Q(\reg_temp[85] ));
 sky130_fd_sc_hd__dfrtp_4 _2166_ (.CLK(clknet_leaf_2_wb_clk_i),
    .D(_0358_),
    .RESET_B(_0101_),
    .Q(\reg_temp[86] ));
 sky130_fd_sc_hd__dfrtp_4 _2167_ (.CLK(clknet_leaf_4_wb_clk_i),
    .D(_0359_),
    .RESET_B(_0102_),
    .Q(\reg_temp[87] ));
 sky130_fd_sc_hd__dfrtp_4 _2168_ (.CLK(clknet_leaf_4_wb_clk_i),
    .D(net1577),
    .RESET_B(_0103_),
    .Q(\reg_temp[88] ));
 sky130_fd_sc_hd__dfrtp_4 _2169_ (.CLK(clknet_leaf_5_wb_clk_i),
    .D(_0361_),
    .RESET_B(_0104_),
    .Q(\reg_temp[89] ));
 sky130_fd_sc_hd__dfrtp_4 _2170_ (.CLK(clknet_leaf_2_wb_clk_i),
    .D(net1552),
    .RESET_B(_0105_),
    .Q(\reg_temp[90] ));
 sky130_fd_sc_hd__dfrtp_4 _2171_ (.CLK(clknet_leaf_0_wb_clk_i),
    .D(net1531),
    .RESET_B(_0106_),
    .Q(\reg_temp[91] ));
 sky130_fd_sc_hd__dfrtp_4 _2172_ (.CLK(clknet_leaf_0_wb_clk_i),
    .D(net1558),
    .RESET_B(_0107_),
    .Q(\reg_temp[92] ));
 sky130_fd_sc_hd__dfrtp_4 _2173_ (.CLK(clknet_leaf_0_wb_clk_i),
    .D(net1536),
    .RESET_B(_0108_),
    .Q(\reg_temp[93] ));
 sky130_fd_sc_hd__dfrtp_4 _2174_ (.CLK(clknet_leaf_2_wb_clk_i),
    .D(net1500),
    .RESET_B(_0109_),
    .Q(\reg_temp[94] ));
 sky130_fd_sc_hd__dfrtp_4 _2175_ (.CLK(clknet_leaf_2_wb_clk_i),
    .D(net1611),
    .RESET_B(_0110_),
    .Q(\reg_temp[95] ));
 sky130_fd_sc_hd__dfrtp_4 _2176_ (.CLK(clknet_leaf_2_wb_clk_i),
    .D(_0368_),
    .RESET_B(_0111_),
    .Q(\reg_temp[96] ));
 sky130_fd_sc_hd__dfrtp_4 _2177_ (.CLK(clknet_leaf_2_wb_clk_i),
    .D(_0369_),
    .RESET_B(_0112_),
    .Q(\reg_temp[97] ));
 sky130_fd_sc_hd__dfrtp_4 _2178_ (.CLK(clknet_leaf_8_wb_clk_i),
    .D(_0370_),
    .RESET_B(_0113_),
    .Q(\reg_temp[98] ));
 sky130_fd_sc_hd__dfrtp_4 _2179_ (.CLK(clknet_leaf_6_wb_clk_i),
    .D(_0371_),
    .RESET_B(_0114_),
    .Q(\reg_temp[99] ));
 sky130_fd_sc_hd__dfrtp_4 _2180_ (.CLK(clknet_leaf_6_wb_clk_i),
    .D(_0372_),
    .RESET_B(_0115_),
    .Q(\reg_temp[100] ));
 sky130_fd_sc_hd__dfrtp_4 _2181_ (.CLK(clknet_leaf_5_wb_clk_i),
    .D(_0373_),
    .RESET_B(_0116_),
    .Q(\reg_temp[101] ));
 sky130_fd_sc_hd__dfrtp_4 _2182_ (.CLK(clknet_leaf_5_wb_clk_i),
    .D(_0374_),
    .RESET_B(_0117_),
    .Q(\reg_temp[102] ));
 sky130_fd_sc_hd__dfrtp_4 _2183_ (.CLK(clknet_leaf_6_wb_clk_i),
    .D(_0375_),
    .RESET_B(_0118_),
    .Q(\reg_temp[103] ));
 sky130_fd_sc_hd__dfrtp_4 _2184_ (.CLK(clknet_leaf_6_wb_clk_i),
    .D(_0376_),
    .RESET_B(_0119_),
    .Q(\reg_temp[104] ));
 sky130_fd_sc_hd__dfrtp_4 _2185_ (.CLK(clknet_leaf_1_wb_clk_i),
    .D(_0377_),
    .RESET_B(_0120_),
    .Q(\reg_temp[105] ));
 sky130_fd_sc_hd__dfrtp_4 _2186_ (.CLK(clknet_leaf_1_wb_clk_i),
    .D(net786),
    .RESET_B(_0121_),
    .Q(\reg_temp[106] ));
 sky130_fd_sc_hd__dfrtp_4 _2187_ (.CLK(clknet_leaf_8_wb_clk_i),
    .D(net869),
    .RESET_B(_0122_),
    .Q(\reg_temp[107] ));
 sky130_fd_sc_hd__dfrtp_4 _2188_ (.CLK(clknet_leaf_8_wb_clk_i),
    .D(net907),
    .RESET_B(_0123_),
    .Q(\reg_temp[108] ));
 sky130_fd_sc_hd__dfrtp_4 _2189_ (.CLK(clknet_leaf_6_wb_clk_i),
    .D(_0381_),
    .RESET_B(_0124_),
    .Q(\reg_temp[109] ));
 sky130_fd_sc_hd__dfrtp_4 _2190_ (.CLK(clknet_leaf_6_wb_clk_i),
    .D(_0382_),
    .RESET_B(_0125_),
    .Q(\reg_temp[110] ));
 sky130_fd_sc_hd__dfrtp_4 _2191_ (.CLK(clknet_leaf_6_wb_clk_i),
    .D(net1573),
    .RESET_B(_0126_),
    .Q(\reg_temp[111] ));
 sky130_fd_sc_hd__dfrtp_4 _2192_ (.CLK(clknet_leaf_6_wb_clk_i),
    .D(_0384_),
    .RESET_B(_0127_),
    .Q(\reg_temp[112] ));
 sky130_fd_sc_hd__dfrtp_4 _2193_ (.CLK(clknet_leaf_7_wb_clk_i),
    .D(_0385_),
    .RESET_B(_0128_),
    .Q(\reg_temp[113] ));
 sky130_fd_sc_hd__dfrtp_4 _2194_ (.CLK(clknet_leaf_6_wb_clk_i),
    .D(net1617),
    .RESET_B(_0129_),
    .Q(\reg_temp[114] ));
 sky130_fd_sc_hd__dfrtp_4 _2195_ (.CLK(clknet_leaf_7_wb_clk_i),
    .D(_0387_),
    .RESET_B(_0130_),
    .Q(\reg_temp[115] ));
 sky130_fd_sc_hd__dfrtp_4 _2196_ (.CLK(clknet_leaf_7_wb_clk_i),
    .D(net1593),
    .RESET_B(_0131_),
    .Q(\reg_temp[116] ));
 sky130_fd_sc_hd__dfrtp_4 _2197_ (.CLK(clknet_leaf_7_wb_clk_i),
    .D(net1570),
    .RESET_B(_0132_),
    .Q(\reg_temp[117] ));
 sky130_fd_sc_hd__dfrtp_4 _2198_ (.CLK(clknet_leaf_8_wb_clk_i),
    .D(net1566),
    .RESET_B(_0133_),
    .Q(\reg_temp[118] ));
 sky130_fd_sc_hd__dfrtp_4 _2199_ (.CLK(clknet_leaf_8_wb_clk_i),
    .D(_0391_),
    .RESET_B(_0134_),
    .Q(\reg_temp[119] ));
 sky130_fd_sc_hd__dfrtp_4 _2200_ (.CLK(clknet_leaf_1_wb_clk_i),
    .D(_0392_),
    .RESET_B(_0135_),
    .Q(\reg_temp[120] ));
 sky130_fd_sc_hd__dfrtp_4 _2201_ (.CLK(clknet_leaf_1_wb_clk_i),
    .D(_0393_),
    .RESET_B(_0136_),
    .Q(\reg_temp[121] ));
 sky130_fd_sc_hd__dfrtp_4 _2202_ (.CLK(clknet_leaf_1_wb_clk_i),
    .D(net1527),
    .RESET_B(_0137_),
    .Q(\reg_temp[122] ));
 sky130_fd_sc_hd__dfrtp_4 _2203_ (.CLK(clknet_leaf_24_wb_clk_i),
    .D(net1549),
    .RESET_B(_0138_),
    .Q(\reg_temp[123] ));
 sky130_fd_sc_hd__dfrtp_4 _2204_ (.CLK(clknet_leaf_23_wb_clk_i),
    .D(net731),
    .RESET_B(_0139_),
    .Q(\reg_temp[124] ));
 sky130_fd_sc_hd__dfrtp_4 _2205_ (.CLK(clknet_leaf_23_wb_clk_i),
    .D(net703),
    .RESET_B(_0140_),
    .Q(\reg_temp[125] ));
 sky130_fd_sc_hd__dfrtp_4 _2206_ (.CLK(clknet_leaf_1_wb_clk_i),
    .D(_0398_),
    .RESET_B(_0141_),
    .Q(\reg_temp[126] ));
 sky130_fd_sc_hd__dfrtp_4 _2207_ (.CLK(clknet_leaf_23_wb_clk_i),
    .D(net671),
    .RESET_B(_0142_),
    .Q(\reg_temp[127] ));
 sky130_fd_sc_hd__dfrtp_4 _2208_ (.CLK(clknet_leaf_23_wb_clk_i),
    .D(net718),
    .RESET_B(_0143_),
    .Q(\reg_temp[128] ));
 sky130_fd_sc_hd__dfrtp_4 _2209_ (.CLK(clknet_leaf_1_wb_clk_i),
    .D(net754),
    .RESET_B(_0144_),
    .Q(\reg_temp[129] ));
 sky130_fd_sc_hd__dfrtp_4 _2210_ (.CLK(clknet_leaf_1_wb_clk_i),
    .D(net800),
    .RESET_B(_0145_),
    .Q(\reg_temp[130] ));
 sky130_fd_sc_hd__dfrtp_2 _2211_ (.CLK(clknet_leaf_9_wb_clk_i),
    .D(net915),
    .RESET_B(_0146_),
    .Q(\reg_temp[131] ));
 sky130_fd_sc_hd__dfrtp_4 _2212_ (.CLK(clknet_leaf_1_wb_clk_i),
    .D(net823),
    .RESET_B(_0147_),
    .Q(\reg_temp[132] ));
 sky130_fd_sc_hd__dfrtp_4 _2213_ (.CLK(clknet_leaf_8_wb_clk_i),
    .D(net925),
    .RESET_B(_0148_),
    .Q(\reg_temp[133] ));
 sky130_fd_sc_hd__dfrtp_4 _2214_ (.CLK(clknet_leaf_8_wb_clk_i),
    .D(net944),
    .RESET_B(_0149_),
    .Q(\reg_temp[134] ));
 sky130_fd_sc_hd__dfrtp_4 _2215_ (.CLK(clknet_leaf_7_wb_clk_i),
    .D(net1012),
    .RESET_B(_0150_),
    .Q(\reg_temp[135] ));
 sky130_fd_sc_hd__dfrtp_2 _2216_ (.CLK(clknet_leaf_7_wb_clk_i),
    .D(net1097),
    .RESET_B(_0151_),
    .Q(\reg_temp[136] ));
 sky130_fd_sc_hd__dfrtp_4 _2217_ (.CLK(clknet_leaf_7_wb_clk_i),
    .D(net1541),
    .RESET_B(_0152_),
    .Q(\reg_temp[137] ));
 sky130_fd_sc_hd__dfrtp_4 _2218_ (.CLK(clknet_leaf_11_wb_clk_i),
    .D(_0410_),
    .RESET_B(_0153_),
    .Q(\reg_temp[138] ));
 sky130_fd_sc_hd__dfrtp_4 _2219_ (.CLK(clknet_leaf_8_wb_clk_i),
    .D(_0411_),
    .RESET_B(_0154_),
    .Q(\reg_temp[139] ));
 sky130_fd_sc_hd__dfrtp_4 _2220_ (.CLK(clknet_leaf_9_wb_clk_i),
    .D(net1140),
    .RESET_B(_0155_),
    .Q(\reg_temp[140] ));
 sky130_fd_sc_hd__dfrtp_4 _2221_ (.CLK(clknet_leaf_10_wb_clk_i),
    .D(net1124),
    .RESET_B(_0156_),
    .Q(\reg_temp[141] ));
 sky130_fd_sc_hd__dfrtp_2 _2222_ (.CLK(clknet_leaf_10_wb_clk_i),
    .D(net1159),
    .RESET_B(_0157_),
    .Q(\reg_temp[142] ));
 sky130_fd_sc_hd__dfrtp_4 _2223_ (.CLK(clknet_leaf_11_wb_clk_i),
    .D(_0415_),
    .RESET_B(_0158_),
    .Q(\reg_temp[143] ));
 sky130_fd_sc_hd__dfrtp_2 _2224_ (.CLK(clknet_leaf_12_wb_clk_i),
    .D(net986),
    .RESET_B(_0159_),
    .Q(\reg_temp[144] ));
 sky130_fd_sc_hd__dfrtp_2 _2225_ (.CLK(clknet_leaf_10_wb_clk_i),
    .D(net1136),
    .RESET_B(_0160_),
    .Q(\reg_temp[145] ));
 sky130_fd_sc_hd__dfrtp_2 _2226_ (.CLK(clknet_leaf_14_wb_clk_i),
    .D(_0418_),
    .RESET_B(_0161_),
    .Q(\reg_temp[146] ));
 sky130_fd_sc_hd__dfrtp_1 _2227_ (.CLK(clknet_leaf_14_wb_clk_i),
    .D(net984),
    .RESET_B(_0162_),
    .Q(\reg_temp[147] ));
 sky130_fd_sc_hd__dfrtp_1 _2228_ (.CLK(clknet_leaf_18_wb_clk_i),
    .D(net971),
    .RESET_B(_0163_),
    .Q(\reg_temp[148] ));
 sky130_fd_sc_hd__dfrtp_1 _2229_ (.CLK(clknet_leaf_18_wb_clk_i),
    .D(net1053),
    .RESET_B(_0164_),
    .Q(\reg_temp[149] ));
 sky130_fd_sc_hd__dfrtp_1 _2230_ (.CLK(clknet_leaf_14_wb_clk_i),
    .D(net1018),
    .RESET_B(_0165_),
    .Q(\reg_temp[150] ));
 sky130_fd_sc_hd__dfrtp_1 _2231_ (.CLK(clknet_leaf_14_wb_clk_i),
    .D(net1112),
    .RESET_B(_0166_),
    .Q(\reg_temp[151] ));
 sky130_fd_sc_hd__dfrtp_1 _2232_ (.CLK(clknet_leaf_14_wb_clk_i),
    .D(net1076),
    .RESET_B(_0167_),
    .Q(\reg_temp[152] ));
 sky130_fd_sc_hd__dfrtp_1 _2233_ (.CLK(clknet_leaf_13_wb_clk_i),
    .D(net1055),
    .RESET_B(_0168_),
    .Q(\reg_temp[153] ));
 sky130_fd_sc_hd__dfrtp_1 _2234_ (.CLK(clknet_leaf_13_wb_clk_i),
    .D(net1020),
    .RESET_B(_0169_),
    .Q(\reg_temp[154] ));
 sky130_fd_sc_hd__dfrtp_1 _2235_ (.CLK(clknet_leaf_13_wb_clk_i),
    .D(net1104),
    .RESET_B(_0170_),
    .Q(\reg_temp[155] ));
 sky130_fd_sc_hd__dfrtp_1 _2236_ (.CLK(clknet_leaf_13_wb_clk_i),
    .D(net1102),
    .RESET_B(_0171_),
    .Q(\reg_temp[156] ));
 sky130_fd_sc_hd__dfrtp_1 _2237_ (.CLK(clknet_leaf_13_wb_clk_i),
    .D(net1175),
    .RESET_B(_0172_),
    .Q(\reg_temp[157] ));
 sky130_fd_sc_hd__dfrtp_1 _2238_ (.CLK(clknet_leaf_13_wb_clk_i),
    .D(net1074),
    .RESET_B(_0173_),
    .Q(\reg_temp[158] ));
 sky130_fd_sc_hd__dfrtp_1 _2239_ (.CLK(clknet_leaf_14_wb_clk_i),
    .D(net961),
    .RESET_B(_0174_),
    .Q(\reg_temp[159] ));
 sky130_fd_sc_hd__dfrtp_1 _2240_ (.CLK(clknet_leaf_18_wb_clk_i),
    .D(net898),
    .RESET_B(_0175_),
    .Q(\reg_temp[160] ));
 sky130_fd_sc_hd__dfrtp_1 _2241_ (.CLK(clknet_leaf_18_wb_clk_i),
    .D(net872),
    .RESET_B(_0176_),
    .Q(\reg_temp[161] ));
 sky130_fd_sc_hd__dfrtp_1 _2242_ (.CLK(clknet_leaf_18_wb_clk_i),
    .D(net930),
    .RESET_B(_0177_),
    .Q(\reg_temp[162] ));
 sky130_fd_sc_hd__dlxtn_1 _2243_ (.D(_0003_),
    .GATE_N(net572),
    .Q(updateRegs));
 sky130_fd_sc_hd__dfrtp_1 _2244_ (.CLK(clknet_leaf_25_wb_clk_i),
    .D(net661),
    .RESET_B(_0178_),
    .Q(net516));
 sky130_fd_sc_hd__dfrtp_1 _2245_ (.CLK(clknet_leaf_25_wb_clk_i),
    .D(net1207),
    .RESET_B(_0179_),
    .Q(net517));
 sky130_fd_sc_hd__dfrtp_1 _2246_ (.CLK(clknet_leaf_25_wb_clk_i),
    .D(net1214),
    .RESET_B(_0180_),
    .Q(net518));
 sky130_fd_sc_hd__dfrtp_2 _2247_ (.CLK(clknet_leaf_25_wb_clk_i),
    .D(net1153),
    .RESET_B(_0181_),
    .Q(net520));
 sky130_fd_sc_hd__dfrtp_4 _2248_ (.CLK(clknet_leaf_25_wb_clk_i),
    .D(\next_state[0] ),
    .RESET_B(_0182_),
    .Q(\current_state[0] ));
 sky130_fd_sc_hd__dfrtp_2 _2249_ (.CLK(clknet_leaf_25_wb_clk_i),
    .D(\next_state[1] ),
    .RESET_B(_0183_),
    .Q(\current_state[1] ));
 sky130_fd_sc_hd__dfrtp_1 _2250_ (.CLK(clknet_leaf_22_wb_clk_i),
    .D(_0439_),
    .RESET_B(_0184_),
    .Q(net447));
 sky130_fd_sc_hd__dfrtp_1 _2251_ (.CLK(clknet_leaf_24_wb_clk_i),
    .D(_0440_),
    .RESET_B(_0185_),
    .Q(net448));
 sky130_fd_sc_hd__dfrtp_1 _2252_ (.CLK(clknet_leaf_22_wb_clk_i),
    .D(_0441_),
    .RESET_B(_0186_),
    .Q(net449));
 sky130_fd_sc_hd__dfrtp_1 _2253_ (.CLK(clknet_leaf_23_wb_clk_i),
    .D(_0442_),
    .RESET_B(_0187_),
    .Q(net450));
 sky130_fd_sc_hd__dfrtp_1 _2254_ (.CLK(clknet_leaf_23_wb_clk_i),
    .D(_0443_),
    .RESET_B(_0188_),
    .Q(net451));
 sky130_fd_sc_hd__dfrtp_1 _2255_ (.CLK(clknet_leaf_22_wb_clk_i),
    .D(_0444_),
    .RESET_B(_0189_),
    .Q(net452));
 sky130_fd_sc_hd__dfrtp_1 _2256_ (.CLK(clknet_leaf_9_wb_clk_i),
    .D(_0445_),
    .RESET_B(_0190_),
    .Q(net453));
 sky130_fd_sc_hd__dfrtp_1 _2257_ (.CLK(clknet_leaf_23_wb_clk_i),
    .D(_0446_),
    .RESET_B(_0191_),
    .Q(net454));
 sky130_fd_sc_hd__dfrtp_1 _2258_ (.CLK(clknet_leaf_16_wb_clk_i),
    .D(_0447_),
    .RESET_B(_0192_),
    .Q(net455));
 sky130_fd_sc_hd__dfrtp_1 _2259_ (.CLK(clknet_leaf_23_wb_clk_i),
    .D(_0448_),
    .RESET_B(_0193_),
    .Q(net456));
 sky130_fd_sc_hd__dfrtp_1 _2260_ (.CLK(clknet_leaf_23_wb_clk_i),
    .D(_0449_),
    .RESET_B(_0194_),
    .Q(net457));
 sky130_fd_sc_hd__dfrtp_1 _2261_ (.CLK(clknet_leaf_23_wb_clk_i),
    .D(_0450_),
    .RESET_B(_0195_),
    .Q(net458));
 sky130_fd_sc_hd__dfrtp_1 _2262_ (.CLK(clknet_leaf_16_wb_clk_i),
    .D(_0451_),
    .RESET_B(_0196_),
    .Q(net459));
 sky130_fd_sc_hd__dfrtp_1 _2263_ (.CLK(clknet_leaf_16_wb_clk_i),
    .D(_0452_),
    .RESET_B(_0197_),
    .Q(net460));
 sky130_fd_sc_hd__dfrtp_1 _2264_ (.CLK(clknet_leaf_22_wb_clk_i),
    .D(net1266),
    .RESET_B(_0198_),
    .Q(net461));
 sky130_fd_sc_hd__dfrtp_1 _2265_ (.CLK(clknet_leaf_22_wb_clk_i),
    .D(_0454_),
    .RESET_B(_0199_),
    .Q(net462));
 sky130_fd_sc_hd__dfrtp_1 _2266_ (.CLK(clknet_leaf_16_wb_clk_i),
    .D(_0455_),
    .RESET_B(_0200_),
    .Q(net463));
 sky130_fd_sc_hd__dfrtp_1 _2267_ (.CLK(clknet_leaf_22_wb_clk_i),
    .D(_0456_),
    .RESET_B(_0201_),
    .Q(net464));
 sky130_fd_sc_hd__dfrtp_1 _2268_ (.CLK(clknet_leaf_15_wb_clk_i),
    .D(_0457_),
    .RESET_B(_0202_),
    .Q(net465));
 sky130_fd_sc_hd__dfrtp_1 _2269_ (.CLK(clknet_leaf_23_wb_clk_i),
    .D(_0458_),
    .RESET_B(_0203_),
    .Q(net466));
 sky130_fd_sc_hd__dfrtp_1 _2270_ (.CLK(clknet_leaf_16_wb_clk_i),
    .D(_0459_),
    .RESET_B(_0204_),
    .Q(net467));
 sky130_fd_sc_hd__dfrtp_1 _2271_ (.CLK(clknet_leaf_22_wb_clk_i),
    .D(_0460_),
    .RESET_B(_0205_),
    .Q(net468));
 sky130_fd_sc_hd__dfrtp_1 _2272_ (.CLK(clknet_leaf_22_wb_clk_i),
    .D(net1222),
    .RESET_B(_0206_),
    .Q(net469));
 sky130_fd_sc_hd__dfrtp_1 _2273_ (.CLK(clknet_leaf_22_wb_clk_i),
    .D(_0462_),
    .RESET_B(_0207_),
    .Q(net470));
 sky130_fd_sc_hd__dfrtp_1 _2274_ (.CLK(clknet_leaf_22_wb_clk_i),
    .D(net1268),
    .RESET_B(_0208_),
    .Q(net471));
 sky130_fd_sc_hd__dfrtp_1 _2275_ (.CLK(clknet_leaf_22_wb_clk_i),
    .D(_0464_),
    .RESET_B(_0209_),
    .Q(net472));
 sky130_fd_sc_hd__dfrtp_1 _2276_ (.CLK(clknet_leaf_22_wb_clk_i),
    .D(net1258),
    .RESET_B(_0210_),
    .Q(net473));
 sky130_fd_sc_hd__dfrtp_1 _2277_ (.CLK(clknet_leaf_22_wb_clk_i),
    .D(_0466_),
    .RESET_B(_0211_),
    .Q(net474));
 sky130_fd_sc_hd__dfrtp_1 _2278_ (.CLK(clknet_leaf_15_wb_clk_i),
    .D(net1226),
    .RESET_B(_0212_),
    .Q(net475));
 sky130_fd_sc_hd__dfrtp_1 _2279_ (.CLK(clknet_leaf_22_wb_clk_i),
    .D(_0468_),
    .RESET_B(_0213_),
    .Q(net476));
 sky130_fd_sc_hd__dfrtp_1 _2280_ (.CLK(clknet_leaf_22_wb_clk_i),
    .D(net1270),
    .RESET_B(_0214_),
    .Q(net477));
 sky130_fd_sc_hd__dfrtp_1 _2281_ (.CLK(clknet_leaf_22_wb_clk_i),
    .D(_0470_),
    .RESET_B(_0215_),
    .Q(net478));
 sky130_fd_sc_hd__dfrtp_1 _2282_ (.CLK(clknet_leaf_16_wb_clk_i),
    .D(_0471_),
    .RESET_B(_0216_),
    .Q(net479));
 sky130_fd_sc_hd__dfrtp_1 _2283_ (.CLK(clknet_leaf_15_wb_clk_i),
    .D(_0472_),
    .RESET_B(_0217_),
    .Q(net480));
 sky130_fd_sc_hd__dfrtp_1 _2284_ (.CLK(clknet_leaf_21_wb_clk_i),
    .D(_0473_),
    .RESET_B(_0218_),
    .Q(net481));
 sky130_fd_sc_hd__dfrtp_1 _2285_ (.CLK(clknet_leaf_21_wb_clk_i),
    .D(_0474_),
    .RESET_B(_0219_),
    .Q(net482));
 sky130_fd_sc_hd__dfrtp_1 _2286_ (.CLK(clknet_leaf_15_wb_clk_i),
    .D(_0475_),
    .RESET_B(_0220_),
    .Q(net483));
 sky130_fd_sc_hd__dfrtp_1 _2287_ (.CLK(clknet_leaf_15_wb_clk_i),
    .D(_0476_),
    .RESET_B(_0221_),
    .Q(net484));
 sky130_fd_sc_hd__dfrtp_1 _2288_ (.CLK(clknet_leaf_16_wb_clk_i),
    .D(_0477_),
    .RESET_B(_0222_),
    .Q(net485));
 sky130_fd_sc_hd__dfrtp_1 _2289_ (.CLK(clknet_leaf_22_wb_clk_i),
    .D(_0478_),
    .RESET_B(_0223_),
    .Q(net486));
 sky130_fd_sc_hd__dfrtp_1 _2290_ (.CLK(clknet_leaf_21_wb_clk_i),
    .D(net1279),
    .RESET_B(_0224_),
    .Q(net487));
 sky130_fd_sc_hd__dfrtp_1 _2291_ (.CLK(clknet_leaf_22_wb_clk_i),
    .D(_0480_),
    .RESET_B(_0225_),
    .Q(net488));
 sky130_fd_sc_hd__dfrtp_1 _2292_ (.CLK(clknet_leaf_21_wb_clk_i),
    .D(_0481_),
    .RESET_B(_0226_),
    .Q(net489));
 sky130_fd_sc_hd__dfrtp_1 _2293_ (.CLK(clknet_leaf_21_wb_clk_i),
    .D(_0482_),
    .RESET_B(_0227_),
    .Q(net490));
 sky130_fd_sc_hd__dfrtp_1 _2294_ (.CLK(clknet_leaf_21_wb_clk_i),
    .D(net1276),
    .RESET_B(_0228_),
    .Q(net491));
 sky130_fd_sc_hd__dfrtp_1 _2295_ (.CLK(clknet_leaf_16_wb_clk_i),
    .D(_0484_),
    .RESET_B(_0229_),
    .Q(net492));
 sky130_fd_sc_hd__dfrtp_1 _2296_ (.CLK(clknet_leaf_16_wb_clk_i),
    .D(_0485_),
    .RESET_B(_0230_),
    .Q(net493));
 sky130_fd_sc_hd__dfrtp_1 _2297_ (.CLK(clknet_leaf_19_wb_clk_i),
    .D(_0486_),
    .RESET_B(_0231_),
    .Q(net494));
 sky130_fd_sc_hd__dfrtp_1 _2298_ (.CLK(clknet_leaf_17_wb_clk_i),
    .D(_0487_),
    .RESET_B(_0232_),
    .Q(net495));
 sky130_fd_sc_hd__dfrtp_1 _2299_ (.CLK(clknet_leaf_17_wb_clk_i),
    .D(_0488_),
    .RESET_B(_0233_),
    .Q(net496));
 sky130_fd_sc_hd__dfrtp_1 _2300_ (.CLK(clknet_leaf_15_wb_clk_i),
    .D(_0489_),
    .RESET_B(_0234_),
    .Q(net497));
 sky130_fd_sc_hd__dfrtp_1 _2301_ (.CLK(clknet_leaf_21_wb_clk_i),
    .D(net1311),
    .RESET_B(_0235_),
    .Q(net498));
 sky130_fd_sc_hd__dfrtp_1 _2302_ (.CLK(clknet_leaf_17_wb_clk_i),
    .D(_0491_),
    .RESET_B(_0236_),
    .Q(net499));
 sky130_fd_sc_hd__dfrtp_1 _2303_ (.CLK(clknet_leaf_21_wb_clk_i),
    .D(net1314),
    .RESET_B(_0237_),
    .Q(net500));
 sky130_fd_sc_hd__dfrtp_1 _2304_ (.CLK(clknet_leaf_20_wb_clk_i),
    .D(net1288),
    .RESET_B(_0238_),
    .Q(net501));
 sky130_fd_sc_hd__dfrtp_1 _2305_ (.CLK(clknet_leaf_20_wb_clk_i),
    .D(_0494_),
    .RESET_B(_0239_),
    .Q(net502));
 sky130_fd_sc_hd__dfrtp_1 _2306_ (.CLK(clknet_leaf_20_wb_clk_i),
    .D(_0495_),
    .RESET_B(_0240_),
    .Q(net503));
 sky130_fd_sc_hd__dfrtp_1 _2307_ (.CLK(clknet_leaf_20_wb_clk_i),
    .D(_0496_),
    .RESET_B(_0241_),
    .Q(net504));
 sky130_fd_sc_hd__dfrtp_1 _2308_ (.CLK(clknet_leaf_19_wb_clk_i),
    .D(_0497_),
    .RESET_B(_0242_),
    .Q(net505));
 sky130_fd_sc_hd__dfrtp_1 _2309_ (.CLK(clknet_leaf_17_wb_clk_i),
    .D(_0498_),
    .RESET_B(_0243_),
    .Q(net506));
 sky130_fd_sc_hd__dfrtp_1 _2310_ (.CLK(clknet_leaf_17_wb_clk_i),
    .D(_0499_),
    .RESET_B(_0244_),
    .Q(net507));
 sky130_fd_sc_hd__dfrtp_1 _2311_ (.CLK(clknet_leaf_20_wb_clk_i),
    .D(net1291),
    .RESET_B(_0245_),
    .Q(net508));
 sky130_fd_sc_hd__dfrtp_1 _2312_ (.CLK(clknet_leaf_21_wb_clk_i),
    .D(_0501_),
    .RESET_B(_0246_),
    .Q(net509));
 sky130_fd_sc_hd__dfrtp_1 _2313_ (.CLK(clknet_leaf_17_wb_clk_i),
    .D(_0502_),
    .RESET_B(_0247_),
    .Q(net510));
 sky130_fd_sc_hd__dfrtp_1 _2314_ (.CLK(clknet_leaf_19_wb_clk_i),
    .D(_0503_),
    .RESET_B(_0248_),
    .Q(net511));
 sky130_fd_sc_hd__dfrtp_1 _2315_ (.CLK(clknet_leaf_17_wb_clk_i),
    .D(_0504_),
    .RESET_B(_0249_),
    .Q(net512));
 sky130_fd_sc_hd__dfrtp_1 _2316_ (.CLK(clknet_leaf_19_wb_clk_i),
    .D(_0505_),
    .RESET_B(_0250_),
    .Q(net513));
 sky130_fd_sc_hd__dfrtp_1 _2317_ (.CLK(clknet_leaf_20_wb_clk_i),
    .D(_0506_),
    .RESET_B(_0251_),
    .Q(net514));
 sky130_fd_sc_hd__dfrtp_1 _2318_ (.CLK(clknet_leaf_20_wb_clk_i),
    .D(_0507_),
    .RESET_B(_0252_),
    .Q(net427));
 sky130_fd_sc_hd__dfrtp_1 _2319_ (.CLK(clknet_leaf_19_wb_clk_i),
    .D(_0508_),
    .RESET_B(_0253_),
    .Q(net428));
 sky130_fd_sc_hd__dfrtp_1 _2320_ (.CLK(clknet_leaf_20_wb_clk_i),
    .D(_0509_),
    .RESET_B(_0254_),
    .Q(net429));
 sky130_fd_sc_hd__dfrtp_1 _2321_ (.CLK(clknet_leaf_19_wb_clk_i),
    .D(_0510_),
    .RESET_B(_0255_),
    .Q(net430));
 sky130_fd_sc_hd__dfrtp_1 _2322_ (.CLK(clknet_leaf_18_wb_clk_i),
    .D(_0511_),
    .RESET_B(_0256_),
    .Q(net431));
 sky130_fd_sc_hd__dfrtp_1 _2323_ (.CLK(clknet_leaf_19_wb_clk_i),
    .D(_0512_),
    .RESET_B(_0257_),
    .Q(net432));
 sky130_fd_sc_hd__dfrtp_1 _2324_ (.CLK(clknet_leaf_19_wb_clk_i),
    .D(_0513_),
    .RESET_B(_0258_),
    .Q(net433));
 sky130_fd_sc_hd__dfrtp_1 _2325_ (.CLK(clknet_leaf_20_wb_clk_i),
    .D(_0514_),
    .RESET_B(_0259_),
    .Q(net434));
 sky130_fd_sc_hd__dfrtp_1 _2326_ (.CLK(clknet_leaf_20_wb_clk_i),
    .D(_0515_),
    .RESET_B(_0260_),
    .Q(net435));
 sky130_fd_sc_hd__dfrtp_1 _2327_ (.CLK(clknet_leaf_20_wb_clk_i),
    .D(_0516_),
    .RESET_B(_0261_),
    .Q(net436));
 sky130_fd_sc_hd__dfrtp_1 _2328_ (.CLK(clknet_leaf_20_wb_clk_i),
    .D(_0517_),
    .RESET_B(_0262_),
    .Q(net437));
 sky130_fd_sc_hd__dfrtp_1 _2329_ (.CLK(clknet_leaf_19_wb_clk_i),
    .D(_0518_),
    .RESET_B(_0263_),
    .Q(net438));
 sky130_fd_sc_hd__dfrtp_1 _2330_ (.CLK(clknet_leaf_19_wb_clk_i),
    .D(_0519_),
    .RESET_B(_0264_),
    .Q(net439));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_0_wb_clk_i (.A(wb_clk_i),
    .X(clknet_0_wb_clk_i));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_0__f_wb_clk_i (.A(clknet_0_wb_clk_i),
    .X(clknet_1_0__leaf_wb_clk_i));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_1__f_wb_clk_i (.A(clknet_0_wb_clk_i),
    .X(clknet_1_1__leaf_wb_clk_i));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_0_wb_clk_i (.A(clknet_1_0__leaf_wb_clk_i),
    .X(clknet_leaf_0_wb_clk_i));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_10_wb_clk_i (.A(clknet_1_1__leaf_wb_clk_i),
    .X(clknet_leaf_10_wb_clk_i));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_11_wb_clk_i (.A(clknet_1_1__leaf_wb_clk_i),
    .X(clknet_leaf_11_wb_clk_i));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_12_wb_clk_i (.A(clknet_1_1__leaf_wb_clk_i),
    .X(clknet_leaf_12_wb_clk_i));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_13_wb_clk_i (.A(clknet_1_1__leaf_wb_clk_i),
    .X(clknet_leaf_13_wb_clk_i));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_14_wb_clk_i (.A(clknet_1_1__leaf_wb_clk_i),
    .X(clknet_leaf_14_wb_clk_i));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_15_wb_clk_i (.A(clknet_1_1__leaf_wb_clk_i),
    .X(clknet_leaf_15_wb_clk_i));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_16_wb_clk_i (.A(clknet_1_1__leaf_wb_clk_i),
    .X(clknet_leaf_16_wb_clk_i));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_17_wb_clk_i (.A(clknet_1_1__leaf_wb_clk_i),
    .X(clknet_leaf_17_wb_clk_i));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_18_wb_clk_i (.A(clknet_1_1__leaf_wb_clk_i),
    .X(clknet_leaf_18_wb_clk_i));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_19_wb_clk_i (.A(clknet_1_1__leaf_wb_clk_i),
    .X(clknet_leaf_19_wb_clk_i));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_1_wb_clk_i (.A(clknet_1_0__leaf_wb_clk_i),
    .X(clknet_leaf_1_wb_clk_i));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_20_wb_clk_i (.A(clknet_1_1__leaf_wb_clk_i),
    .X(clknet_leaf_20_wb_clk_i));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_21_wb_clk_i (.A(clknet_1_1__leaf_wb_clk_i),
    .X(clknet_leaf_21_wb_clk_i));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_22_wb_clk_i (.A(clknet_1_1__leaf_wb_clk_i),
    .X(clknet_leaf_22_wb_clk_i));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_23_wb_clk_i (.A(clknet_1_1__leaf_wb_clk_i),
    .X(clknet_leaf_23_wb_clk_i));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_24_wb_clk_i (.A(clknet_1_0__leaf_wb_clk_i),
    .X(clknet_leaf_24_wb_clk_i));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_25_wb_clk_i (.A(clknet_1_0__leaf_wb_clk_i),
    .X(clknet_leaf_25_wb_clk_i));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_26_wb_clk_i (.A(clknet_1_0__leaf_wb_clk_i),
    .X(clknet_leaf_26_wb_clk_i));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_2_wb_clk_i (.A(clknet_1_0__leaf_wb_clk_i),
    .X(clknet_leaf_2_wb_clk_i));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_3_wb_clk_i (.A(clknet_1_0__leaf_wb_clk_i),
    .X(clknet_leaf_3_wb_clk_i));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_4_wb_clk_i (.A(clknet_1_0__leaf_wb_clk_i),
    .X(clknet_leaf_4_wb_clk_i));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_5_wb_clk_i (.A(clknet_1_0__leaf_wb_clk_i),
    .X(clknet_leaf_5_wb_clk_i));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_6_wb_clk_i (.A(clknet_1_0__leaf_wb_clk_i),
    .X(clknet_leaf_6_wb_clk_i));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_7_wb_clk_i (.A(clknet_1_0__leaf_wb_clk_i),
    .X(clknet_leaf_7_wb_clk_i));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_8_wb_clk_i (.A(clknet_1_0__leaf_wb_clk_i),
    .X(clknet_leaf_8_wb_clk_i));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_9_wb_clk_i (.A(clknet_1_0__leaf_wb_clk_i),
    .X(clknet_leaf_9_wb_clk_i));
 sky130_fd_sc_hd__conb_1 controller_618 (.LO(net618));
 sky130_fd_sc_hd__conb_1 controller_619 (.LO(net619));
 sky130_fd_sc_hd__conb_1 controller_620 (.LO(net620));
 sky130_fd_sc_hd__conb_1 controller_621 (.LO(net621));
 sky130_fd_sc_hd__conb_1 controller_622 (.LO(net622));
 sky130_fd_sc_hd__conb_1 controller_623 (.LO(net623));
 sky130_fd_sc_hd__conb_1 controller_624 (.LO(net624));
 sky130_fd_sc_hd__conb_1 controller_625 (.LO(net625));
 sky130_fd_sc_hd__conb_1 controller_626 (.LO(net626));
 sky130_fd_sc_hd__conb_1 controller_627 (.LO(net627));
 sky130_fd_sc_hd__conb_1 controller_628 (.LO(net628));
 sky130_fd_sc_hd__conb_1 controller_629 (.LO(net629));
 sky130_fd_sc_hd__conb_1 controller_630 (.LO(net630));
 sky130_fd_sc_hd__conb_1 controller_631 (.LO(net631));
 sky130_fd_sc_hd__conb_1 controller_632 (.LO(net632));
 sky130_fd_sc_hd__conb_1 controller_633 (.LO(net633));
 sky130_fd_sc_hd__conb_1 controller_634 (.LO(net634));
 sky130_fd_sc_hd__conb_1 controller_635 (.LO(net635));
 sky130_fd_sc_hd__conb_1 controller_636 (.LO(net636));
 sky130_fd_sc_hd__conb_1 controller_637 (.LO(net637));
 sky130_fd_sc_hd__conb_1 controller_638 (.LO(net638));
 sky130_fd_sc_hd__conb_1 controller_639 (.LO(net639));
 sky130_fd_sc_hd__conb_1 controller_640 (.LO(net640));
 sky130_fd_sc_hd__conb_1 controller_641 (.LO(net641));
 sky130_fd_sc_hd__conb_1 controller_642 (.LO(net642));
 sky130_fd_sc_hd__conb_1 controller_643 (.LO(net643));
 sky130_fd_sc_hd__conb_1 controller_644 (.LO(net644));
 sky130_fd_sc_hd__conb_1 controller_645 (.LO(net645));
 sky130_fd_sc_hd__conb_1 controller_646 (.LO(net646));
 sky130_fd_sc_hd__conb_1 controller_647 (.LO(net647));
 sky130_fd_sc_hd__conb_1 controller_648 (.LO(net648));
 sky130_fd_sc_hd__conb_1 controller_649 (.LO(net649));
 sky130_fd_sc_hd__conb_1 controller_650 (.LO(net650));
 sky130_fd_sc_hd__conb_1 controller_651 (.LO(net651));
 sky130_fd_sc_hd__conb_1 controller_652 (.LO(net652));
 sky130_fd_sc_hd__conb_1 controller_653 (.LO(net653));
 sky130_fd_sc_hd__conb_1 controller_654 (.LO(net654));
 sky130_fd_sc_hd__conb_1 controller_655 (.LO(net655));
 sky130_fd_sc_hd__conb_1 controller_656 (.LO(net656));
 sky130_fd_sc_hd__conb_1 controller_657 (.LO(net657));
 sky130_fd_sc_hd__clkbuf_1 fanout521 (.A(net683),
    .X(net521));
 sky130_fd_sc_hd__buf_6 fanout522 (.A(net683),
    .X(net522));
 sky130_fd_sc_hd__clkbuf_4 fanout523 (.A(net683),
    .X(net523));
 sky130_fd_sc_hd__clkbuf_8 fanout524 (.A(net683),
    .X(net524));
 sky130_fd_sc_hd__buf_6 fanout525 (.A(net683),
    .X(net525));
 sky130_fd_sc_hd__buf_6 fanout526 (.A(net697),
    .X(net526));
 sky130_fd_sc_hd__buf_4 fanout527 (.A(net530),
    .X(net527));
 sky130_fd_sc_hd__buf_2 fanout528 (.A(net530),
    .X(net528));
 sky130_fd_sc_hd__buf_4 fanout529 (.A(net530),
    .X(net529));
 sky130_fd_sc_hd__clkbuf_4 fanout530 (.A(_0588_),
    .X(net530));
 sky130_fd_sc_hd__buf_4 fanout531 (.A(net533),
    .X(net531));
 sky130_fd_sc_hd__clkbuf_4 fanout532 (.A(net533),
    .X(net532));
 sky130_fd_sc_hd__clkbuf_4 fanout533 (.A(_0588_),
    .X(net533));
 sky130_fd_sc_hd__clkbuf_8 fanout534 (.A(net737),
    .X(net534));
 sky130_fd_sc_hd__clkbuf_8 fanout535 (.A(net738),
    .X(net535));
 sky130_fd_sc_hd__clkbuf_1 fanout536 (.A(net737),
    .X(net536));
 sky130_fd_sc_hd__clkbuf_2 fanout537 (.A(net736),
    .X(net537));
 sky130_fd_sc_hd__buf_6 fanout538 (.A(net539),
    .X(net538));
 sky130_fd_sc_hd__clkbuf_8 fanout539 (.A(net736),
    .X(net539));
 sky130_fd_sc_hd__clkbuf_4 fanout540 (.A(net544),
    .X(net540));
 sky130_fd_sc_hd__clkbuf_4 fanout541 (.A(net542),
    .X(net541));
 sky130_fd_sc_hd__clkbuf_4 fanout542 (.A(net544),
    .X(net542));
 sky130_fd_sc_hd__clkbuf_4 fanout543 (.A(net544),
    .X(net543));
 sky130_fd_sc_hd__clkbuf_4 fanout544 (.A(_0946_),
    .X(net544));
 sky130_fd_sc_hd__clkbuf_4 fanout545 (.A(net546),
    .X(net545));
 sky130_fd_sc_hd__clkbuf_4 fanout546 (.A(net551),
    .X(net546));
 sky130_fd_sc_hd__clkbuf_4 fanout547 (.A(net548),
    .X(net547));
 sky130_fd_sc_hd__clkbuf_4 fanout548 (.A(net551),
    .X(net548));
 sky130_fd_sc_hd__clkbuf_4 fanout549 (.A(net550),
    .X(net549));
 sky130_fd_sc_hd__clkbuf_4 fanout550 (.A(net551),
    .X(net550));
 sky130_fd_sc_hd__clkbuf_4 fanout551 (.A(_0946_),
    .X(net551));
 sky130_fd_sc_hd__buf_4 fanout552 (.A(net555),
    .X(net552));
 sky130_fd_sc_hd__clkbuf_4 fanout553 (.A(net555),
    .X(net553));
 sky130_fd_sc_hd__buf_4 fanout554 (.A(net555),
    .X(net554));
 sky130_fd_sc_hd__clkbuf_4 fanout555 (.A(_0589_),
    .X(net555));
 sky130_fd_sc_hd__buf_4 fanout556 (.A(net558),
    .X(net556));
 sky130_fd_sc_hd__clkbuf_4 fanout557 (.A(net558),
    .X(net557));
 sky130_fd_sc_hd__clkbuf_4 fanout558 (.A(_0589_),
    .X(net558));
 sky130_fd_sc_hd__buf_4 fanout559 (.A(_0569_),
    .X(net559));
 sky130_fd_sc_hd__clkbuf_4 fanout560 (.A(_0569_),
    .X(net560));
 sky130_fd_sc_hd__buf_4 fanout561 (.A(net563),
    .X(net561));
 sky130_fd_sc_hd__clkbuf_4 fanout562 (.A(net563),
    .X(net562));
 sky130_fd_sc_hd__clkbuf_8 fanout563 (.A(_0569_),
    .X(net563));
 sky130_fd_sc_hd__buf_4 fanout564 (.A(net567),
    .X(net564));
 sky130_fd_sc_hd__buf_4 fanout565 (.A(net566),
    .X(net565));
 sky130_fd_sc_hd__buf_4 fanout566 (.A(net567),
    .X(net566));
 sky130_fd_sc_hd__buf_4 fanout567 (.A(_0569_),
    .X(net567));
 sky130_fd_sc_hd__clkbuf_8 fanout568 (.A(net570),
    .X(net568));
 sky130_fd_sc_hd__buf_2 fanout569 (.A(net570),
    .X(net569));
 sky130_fd_sc_hd__clkbuf_4 fanout570 (.A(net571),
    .X(net570));
 sky130_fd_sc_hd__buf_4 fanout571 (.A(_0569_),
    .X(net571));
 sky130_fd_sc_hd__buf_4 fanout572 (.A(_0007_),
    .X(net572));
 sky130_fd_sc_hd__clkbuf_4 fanout573 (.A(_0007_),
    .X(net573));
 sky130_fd_sc_hd__buf_4 fanout574 (.A(net576),
    .X(net574));
 sky130_fd_sc_hd__clkbuf_4 fanout575 (.A(net576),
    .X(net575));
 sky130_fd_sc_hd__clkbuf_8 fanout576 (.A(_0007_),
    .X(net576));
 sky130_fd_sc_hd__buf_4 fanout577 (.A(net580),
    .X(net577));
 sky130_fd_sc_hd__buf_4 fanout578 (.A(net579),
    .X(net578));
 sky130_fd_sc_hd__clkbuf_8 fanout579 (.A(net580),
    .X(net579));
 sky130_fd_sc_hd__clkbuf_4 fanout580 (.A(_0007_),
    .X(net580));
 sky130_fd_sc_hd__clkbuf_8 fanout581 (.A(net583),
    .X(net581));
 sky130_fd_sc_hd__buf_2 fanout582 (.A(net583),
    .X(net582));
 sky130_fd_sc_hd__clkbuf_4 fanout583 (.A(net584),
    .X(net583));
 sky130_fd_sc_hd__buf_4 fanout584 (.A(_0007_),
    .X(net584));
 sky130_fd_sc_hd__clkbuf_8 fanout585 (.A(net588),
    .X(net585));
 sky130_fd_sc_hd__clkbuf_8 fanout586 (.A(net588),
    .X(net586));
 sky130_fd_sc_hd__buf_4 fanout587 (.A(net588),
    .X(net587));
 sky130_fd_sc_hd__buf_4 fanout588 (.A(_0592_),
    .X(net588));
 sky130_fd_sc_hd__clkbuf_8 fanout589 (.A(net590),
    .X(net589));
 sky130_fd_sc_hd__buf_6 fanout590 (.A(_0592_),
    .X(net590));
 sky130_fd_sc_hd__buf_4 fanout591 (.A(net594),
    .X(net591));
 sky130_fd_sc_hd__clkbuf_4 fanout592 (.A(net594),
    .X(net592));
 sky130_fd_sc_hd__clkbuf_2 fanout593 (.A(net594),
    .X(net593));
 sky130_fd_sc_hd__buf_2 fanout594 (.A(_0004_),
    .X(net594));
 sky130_fd_sc_hd__buf_2 fanout595 (.A(net597),
    .X(net595));
 sky130_fd_sc_hd__clkbuf_2 fanout596 (.A(net597),
    .X(net596));
 sky130_fd_sc_hd__buf_4 fanout597 (.A(_0004_),
    .X(net597));
 sky130_fd_sc_hd__buf_8 fanout598 (.A(net599),
    .X(net598));
 sky130_fd_sc_hd__clkbuf_8 fanout599 (.A(net262),
    .X(net599));
 sky130_fd_sc_hd__buf_8 fanout600 (.A(net602),
    .X(net600));
 sky130_fd_sc_hd__buf_8 fanout601 (.A(net602),
    .X(net601));
 sky130_fd_sc_hd__buf_8 fanout602 (.A(net262),
    .X(net602));
 sky130_fd_sc_hd__buf_8 fanout603 (.A(net605),
    .X(net603));
 sky130_fd_sc_hd__buf_8 fanout604 (.A(net605),
    .X(net604));
 sky130_fd_sc_hd__buf_4 fanout605 (.A(net606),
    .X(net605));
 sky130_fd_sc_hd__buf_8 fanout606 (.A(net262),
    .X(net606));
 sky130_fd_sc_hd__buf_8 fanout607 (.A(net609),
    .X(net607));
 sky130_fd_sc_hd__buf_8 fanout608 (.A(net609),
    .X(net608));
 sky130_fd_sc_hd__clkbuf_8 fanout609 (.A(net611),
    .X(net609));
 sky130_fd_sc_hd__buf_8 fanout610 (.A(net611),
    .X(net610));
 sky130_fd_sc_hd__buf_4 fanout611 (.A(net262),
    .X(net611));
 sky130_fd_sc_hd__buf_8 fanout612 (.A(net615),
    .X(net612));
 sky130_fd_sc_hd__buf_8 fanout613 (.A(net615),
    .X(net613));
 sky130_fd_sc_hd__buf_4 fanout614 (.A(net615),
    .X(net614));
 sky130_fd_sc_hd__clkbuf_8 fanout615 (.A(net262),
    .X(net615));
 sky130_fd_sc_hd__buf_8 fanout616 (.A(net617),
    .X(net616));
 sky130_fd_sc_hd__clkbuf_8 fanout617 (.A(net262),
    .X(net617));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1 (.A(net1114),
    .X(net658));
 sky130_fd_sc_hd__dlygate4sd3_1 hold10 (.A(la_data_in[45]),
    .X(net667));
 sky130_fd_sc_hd__dlygate4sd3_1 hold100 (.A(net259),
    .X(net757));
 sky130_fd_sc_hd__buf_1 hold101 (.A(_0826_),
    .X(net758));
 sky130_fd_sc_hd__dlygate4sd3_1 hold102 (.A(_0932_),
    .X(net759));
 sky130_fd_sc_hd__dlygate4sd3_1 hold103 (.A(_0274_),
    .X(net760));
 sky130_fd_sc_hd__dlygate4sd3_1 hold104 (.A(net801),
    .X(net761));
 sky130_fd_sc_hd__dlygate4sd3_1 hold105 (.A(net190),
    .X(net762));
 sky130_fd_sc_hd__dlymetal6s2s_1 hold106 (.A(_0778_),
    .X(net763));
 sky130_fd_sc_hd__dlygate4sd3_1 hold107 (.A(_0779_),
    .X(net764));
 sky130_fd_sc_hd__dlygate4sd3_1 hold108 (.A(la_data_in[94]),
    .X(net765));
 sky130_fd_sc_hd__clkbuf_2 hold109 (.A(net257),
    .X(net766));
 sky130_fd_sc_hd__dlygate4sd3_1 hold11 (.A(net203),
    .X(net668));
 sky130_fd_sc_hd__dlygate4sd3_1 hold110 (.A(_0568_),
    .X(net767));
 sky130_fd_sc_hd__clkdlybuf4s25_1 hold111 (.A(_0854_),
    .X(net768));
 sky130_fd_sc_hd__dlygate4sd3_1 hold112 (.A(_0858_),
    .X(net769));
 sky130_fd_sc_hd__buf_1 hold113 (.A(net736),
    .X(net770));
 sky130_fd_sc_hd__dlygate4sd3_1 hold114 (.A(_0310_),
    .X(net771));
 sky130_fd_sc_hd__dlygate4sd3_1 hold115 (.A(net806),
    .X(net772));
 sky130_fd_sc_hd__dlygate4sd3_1 hold116 (.A(net241),
    .X(net773));
 sky130_fd_sc_hd__dlymetal6s2s_1 hold117 (.A(_0830_),
    .X(net774));
 sky130_fd_sc_hd__dlygate4sd3_1 hold118 (.A(_0831_),
    .X(net775));
 sky130_fd_sc_hd__dlygate4sd3_1 hold119 (.A(net1164),
    .X(net776));
 sky130_fd_sc_hd__dlygate4sd3_1 hold12 (.A(_0754_),
    .X(net669));
 sky130_fd_sc_hd__dlygate4sd3_1 hold120 (.A(net172),
    .X(net777));
 sky130_fd_sc_hd__dlygate4sd3_1 hold121 (.A(_0591_),
    .X(net778));
 sky130_fd_sc_hd__clkdlybuf4s25_1 hold122 (.A(_0593_),
    .X(net779));
 sky130_fd_sc_hd__dlygate4sd3_1 hold123 (.A(_0855_),
    .X(net780));
 sky130_fd_sc_hd__dlygate4sd3_1 hold124 (.A(_0350_),
    .X(net781));
 sky130_fd_sc_hd__dlygate4sd3_1 hold125 (.A(net850),
    .X(net782));
 sky130_fd_sc_hd__dlygate4sd3_1 hold126 (.A(net180),
    .X(net783));
 sky130_fd_sc_hd__dlymetal6s2s_1 hold127 (.A(_0796_),
    .X(net784));
 sky130_fd_sc_hd__dlygate4sd3_1 hold128 (.A(_0797_),
    .X(net785));
 sky130_fd_sc_hd__dlygate4sd3_1 hold129 (.A(_0378_),
    .X(net786));
 sky130_fd_sc_hd__dlygate4sd3_1 hold13 (.A(_0755_),
    .X(net670));
 sky130_fd_sc_hd__dlygate4sd3_1 hold130 (.A(net795),
    .X(net787));
 sky130_fd_sc_hd__dlygate4sd3_1 hold131 (.A(net170),
    .X(net788));
 sky130_fd_sc_hd__dlymetal6s2s_1 hold132 (.A(_0814_),
    .X(net789));
 sky130_fd_sc_hd__dlygate4sd3_1 hold133 (.A(_0815_),
    .X(net790));
 sky130_fd_sc_hd__dlygate4sd3_1 hold134 (.A(net810),
    .X(net791));
 sky130_fd_sc_hd__dlygate4sd3_1 hold135 (.A(net191),
    .X(net792));
 sky130_fd_sc_hd__dlymetal6s2s_1 hold136 (.A(_0776_),
    .X(net793));
 sky130_fd_sc_hd__dlygate4sd3_1 hold137 (.A(_0907_),
    .X(net794));
 sky130_fd_sc_hd__dlygate4sd3_1 hold138 (.A(la_data_in[15]),
    .X(net795));
 sky130_fd_sc_hd__dlygate4sd3_1 hold139 (.A(net808),
    .X(net796));
 sky130_fd_sc_hd__dlygate4sd3_1 hold14 (.A(_0399_),
    .X(net671));
 sky130_fd_sc_hd__dlygate4sd3_1 hold140 (.A(net206),
    .X(net797));
 sky130_fd_sc_hd__buf_1 hold141 (.A(_0748_),
    .X(net798));
 sky130_fd_sc_hd__dlygate4sd3_1 hold142 (.A(_0749_),
    .X(net799));
 sky130_fd_sc_hd__dlygate4sd3_1 hold143 (.A(_0402_),
    .X(net800));
 sky130_fd_sc_hd__dlygate4sd3_1 hold144 (.A(la_data_in[33]),
    .X(net801));
 sky130_fd_sc_hd__dlygate4sd3_1 hold145 (.A(net914),
    .X(net802));
 sky130_fd_sc_hd__dlygate4sd3_1 hold146 (.A(net207),
    .X(net803));
 sky130_fd_sc_hd__buf_1 hold147 (.A(_0746_),
    .X(net804));
 sky130_fd_sc_hd__dlygate4sd3_1 hold148 (.A(_0892_),
    .X(net805));
 sky130_fd_sc_hd__dlygate4sd3_1 hold149 (.A(net1574),
    .X(net806));
 sky130_fd_sc_hd__dlygate4sd3_1 hold15 (.A(net1461),
    .X(net672));
 sky130_fd_sc_hd__dlygate4sd3_1 hold150 (.A(net1497),
    .X(net807));
 sky130_fd_sc_hd__dlygate4sd3_1 hold151 (.A(la_data_in[48]),
    .X(net808));
 sky130_fd_sc_hd__dlygate4sd3_1 hold152 (.A(_0313_),
    .X(net809));
 sky130_fd_sc_hd__dlygate4sd3_1 hold153 (.A(la_data_in[34]),
    .X(net810));
 sky130_fd_sc_hd__dlygate4sd3_1 hold154 (.A(net873),
    .X(net811));
 sky130_fd_sc_hd__dlygate4sd3_1 hold155 (.A(net166),
    .X(net812));
 sky130_fd_sc_hd__buf_1 hold156 (.A(_0822_),
    .X(net813));
 sky130_fd_sc_hd__dlygate4sd3_1 hold157 (.A(_0930_),
    .X(net814));
 sky130_fd_sc_hd__dlygate4sd3_1 hold158 (.A(_0276_),
    .X(net815));
 sky130_fd_sc_hd__dlygate4sd3_1 hold159 (.A(net1501),
    .X(net816));
 sky130_fd_sc_hd__dlygate4sd3_1 hold16 (.A(net186),
    .X(net673));
 sky130_fd_sc_hd__dlygate4sd3_1 hold160 (.A(la_data_in[47]),
    .X(net817));
 sky130_fd_sc_hd__dlygate4sd3_1 hold161 (.A(_0312_),
    .X(net818));
 sky130_fd_sc_hd__dlygate4sd3_1 hold162 (.A(net835),
    .X(net819));
 sky130_fd_sc_hd__dlygate4sd3_1 hold163 (.A(net209),
    .X(net820));
 sky130_fd_sc_hd__buf_1 hold164 (.A(_0744_),
    .X(net821));
 sky130_fd_sc_hd__dlygate4sd3_1 hold165 (.A(_0745_),
    .X(net822));
 sky130_fd_sc_hd__dlygate4sd3_1 hold166 (.A(_0404_),
    .X(net823));
 sky130_fd_sc_hd__dlygate4sd3_1 hold167 (.A(net871),
    .X(net824));
 sky130_fd_sc_hd__dlygate4sd3_1 hold168 (.A(net240),
    .X(net825));
 sky130_fd_sc_hd__buf_1 hold169 (.A(_0686_),
    .X(net826));
 sky130_fd_sc_hd__buf_1 hold17 (.A(_0840_),
    .X(net674));
 sky130_fd_sc_hd__dlygate4sd3_1 hold170 (.A(_0862_),
    .X(net827));
 sky130_fd_sc_hd__dlygate4sd3_1 hold171 (.A(_0344_),
    .X(net828));
 sky130_fd_sc_hd__dlygate4sd3_1 hold172 (.A(net1530),
    .X(net829));
 sky130_fd_sc_hd__dlygate4sd3_1 hold173 (.A(net1557),
    .X(net830));
 sky130_fd_sc_hd__dlygate4sd3_1 hold174 (.A(net870),
    .X(net831));
 sky130_fd_sc_hd__dlygate4sd3_1 hold175 (.A(net197),
    .X(net832));
 sky130_fd_sc_hd__buf_1 hold176 (.A(_0838_),
    .X(net833));
 sky130_fd_sc_hd__dlygate4sd3_1 hold177 (.A(_0938_),
    .X(net834));
 sky130_fd_sc_hd__dlygate4sd3_1 hold178 (.A(la_data_in[50]),
    .X(net835));
 sky130_fd_sc_hd__dlygate4sd3_1 hold179 (.A(_0315_),
    .X(net836));
 sky130_fd_sc_hd__dlygate4sd3_1 hold18 (.A(_0939_),
    .X(net675));
 sky130_fd_sc_hd__dlygate4sd3_1 hold180 (.A(net1538),
    .X(net837));
 sky130_fd_sc_hd__dlygate4sd3_1 hold181 (.A(net867),
    .X(net838));
 sky130_fd_sc_hd__dlygate4sd3_1 hold182 (.A(net199),
    .X(net839));
 sky130_fd_sc_hd__buf_1 hold183 (.A(_0762_),
    .X(net840));
 sky130_fd_sc_hd__dlygate4sd3_1 hold184 (.A(_0900_),
    .X(net841));
 sky130_fd_sc_hd__dlygate4sd3_1 hold185 (.A(net862),
    .X(net842));
 sky130_fd_sc_hd__dlygate4sd3_1 hold186 (.A(net252),
    .X(net843));
 sky130_fd_sc_hd__buf_1 hold187 (.A(_0828_),
    .X(net844));
 sky130_fd_sc_hd__dlygate4sd3_1 hold188 (.A(_0933_),
    .X(net845));
 sky130_fd_sc_hd__dlygate4sd3_1 hold189 (.A(net851),
    .X(net846));
 sky130_fd_sc_hd__dlygate4sd3_1 hold19 (.A(_0267_),
    .X(net676));
 sky130_fd_sc_hd__dlygate4sd3_1 hold190 (.A(net198),
    .X(net847));
 sky130_fd_sc_hd__buf_1 hold191 (.A(_0764_),
    .X(net848));
 sky130_fd_sc_hd__dlygate4sd3_1 hold192 (.A(_0901_),
    .X(net849));
 sky130_fd_sc_hd__dlygate4sd3_1 hold193 (.A(la_data_in[24]),
    .X(net850));
 sky130_fd_sc_hd__dlygate4sd3_1 hold194 (.A(net1526),
    .X(net851));
 sky130_fd_sc_hd__dlygate4sd3_1 hold195 (.A(net916),
    .X(net852));
 sky130_fd_sc_hd__dlygate4sd3_1 hold196 (.A(net202),
    .X(net853));
 sky130_fd_sc_hd__buf_1 hold197 (.A(_0756_),
    .X(net854));
 sky130_fd_sc_hd__dlygate4sd3_1 hold198 (.A(_0757_),
    .X(net855));
 sky130_fd_sc_hd__dlygate4sd3_1 hold199 (.A(la_data_in[46]),
    .X(net856));
 sky130_fd_sc_hd__clkbuf_2 hold2 (.A(net174),
    .X(net659));
 sky130_fd_sc_hd__dlygate4sd3_1 hold20 (.A(la_data_in[95]),
    .X(net677));
 sky130_fd_sc_hd__dlygate4sd3_1 hold200 (.A(_0311_),
    .X(net857));
 sky130_fd_sc_hd__dlygate4sd3_1 hold201 (.A(net896),
    .X(net858));
 sky130_fd_sc_hd__dlygate4sd3_1 hold202 (.A(net167),
    .X(net859));
 sky130_fd_sc_hd__buf_1 hold203 (.A(_0820_),
    .X(net860));
 sky130_fd_sc_hd__dlygate4sd3_1 hold204 (.A(_0929_),
    .X(net861));
 sky130_fd_sc_hd__dlygate4sd3_1 hold205 (.A(net1551),
    .X(net862));
 sky130_fd_sc_hd__dlygate4sd3_1 hold206 (.A(net868),
    .X(net863));
 sky130_fd_sc_hd__dlygate4sd3_1 hold207 (.A(net181),
    .X(net864));
 sky130_fd_sc_hd__dlymetal6s2s_1 hold208 (.A(_0794_),
    .X(net865));
 sky130_fd_sc_hd__dlygate4sd3_1 hold209 (.A(_0916_),
    .X(net866));
 sky130_fd_sc_hd__clkbuf_2 hold21 (.A(net258),
    .X(net678));
 sky130_fd_sc_hd__dlygate4sd3_1 hold210 (.A(net1548),
    .X(net867));
 sky130_fd_sc_hd__dlygate4sd3_1 hold211 (.A(la_data_in[25]),
    .X(net868));
 sky130_fd_sc_hd__dlygate4sd3_1 hold212 (.A(_0379_),
    .X(net869));
 sky130_fd_sc_hd__dlygate4sd3_1 hold213 (.A(net1555),
    .X(net870));
 sky130_fd_sc_hd__dlygate4sd3_1 hold214 (.A(la_data_in[79]),
    .X(net871));
 sky130_fd_sc_hd__dlygate4sd3_1 hold215 (.A(_0433_),
    .X(net872));
 sky130_fd_sc_hd__dlygate4sd3_1 hold216 (.A(net1535),
    .X(net873));
 sky130_fd_sc_hd__dlygate4sd3_1 hold217 (.A(net891),
    .X(net874));
 sky130_fd_sc_hd__dlygate4sd3_1 hold218 (.A(net168),
    .X(net875));
 sky130_fd_sc_hd__buf_1 hold219 (.A(_0818_),
    .X(net876));
 sky130_fd_sc_hd__buf_1 hold22 (.A(_0565_),
    .X(net679));
 sky130_fd_sc_hd__dlygate4sd3_1 hold220 (.A(_0928_),
    .X(net877));
 sky130_fd_sc_hd__dlygate4sd3_1 hold221 (.A(net913),
    .X(net878));
 sky130_fd_sc_hd__dlygate4sd3_1 hold222 (.A(net184),
    .X(net879));
 sky130_fd_sc_hd__dlymetal6s2s_1 hold223 (.A(_0788_),
    .X(net880));
 sky130_fd_sc_hd__dlygate4sd3_1 hold224 (.A(_0913_),
    .X(net881));
 sky130_fd_sc_hd__dlygate4sd3_1 hold225 (.A(net959),
    .X(net882));
 sky130_fd_sc_hd__dlygate4sd3_1 hold226 (.A(net195),
    .X(net883));
 sky130_fd_sc_hd__buf_1 hold227 (.A(_0768_),
    .X(net884));
 sky130_fd_sc_hd__dlygate4sd3_1 hold228 (.A(_0769_),
    .X(net885));
 sky130_fd_sc_hd__dlygate4sd3_1 hold229 (.A(net897),
    .X(net886));
 sky130_fd_sc_hd__dlygate4sd3_1 hold23 (.A(_0566_),
    .X(net680));
 sky130_fd_sc_hd__dlygate4sd3_1 hold230 (.A(net239),
    .X(net887));
 sky130_fd_sc_hd__buf_1 hold231 (.A(_0688_),
    .X(net888));
 sky130_fd_sc_hd__dlygate4sd3_1 hold232 (.A(_0863_),
    .X(net889));
 sky130_fd_sc_hd__dlygate4sd3_1 hold233 (.A(_0343_),
    .X(net890));
 sky130_fd_sc_hd__dlygate4sd3_1 hold234 (.A(la_data_in[13]),
    .X(net891));
 sky130_fd_sc_hd__dlygate4sd3_1 hold235 (.A(net919),
    .X(net892));
 sky130_fd_sc_hd__dlygate4sd3_1 hold236 (.A(net183),
    .X(net893));
 sky130_fd_sc_hd__dlymetal6s2s_1 hold237 (.A(_0790_),
    .X(net894));
 sky130_fd_sc_hd__dlygate4sd3_1 hold238 (.A(_0914_),
    .X(net895));
 sky130_fd_sc_hd__dlygate4sd3_1 hold239 (.A(net1499),
    .X(net896));
 sky130_fd_sc_hd__dlygate4sd3_1 hold24 (.A(_0682_),
    .X(net681));
 sky130_fd_sc_hd__dlygate4sd3_1 hold240 (.A(la_data_in[78]),
    .X(net897));
 sky130_fd_sc_hd__dlygate4sd3_1 hold241 (.A(_0432_),
    .X(net898));
 sky130_fd_sc_hd__dlygate4sd3_1 hold242 (.A(net917),
    .X(net899));
 sky130_fd_sc_hd__dlygate4sd3_1 hold243 (.A(net188),
    .X(net900));
 sky130_fd_sc_hd__dlymetal6s2s_1 hold244 (.A(_0782_),
    .X(net901));
 sky130_fd_sc_hd__dlygate4sd3_1 hold245 (.A(_0910_),
    .X(net902));
 sky130_fd_sc_hd__dlygate4sd3_1 hold246 (.A(net908),
    .X(net903));
 sky130_fd_sc_hd__dlygate4sd3_1 hold247 (.A(net182),
    .X(net904));
 sky130_fd_sc_hd__dlymetal6s2s_1 hold248 (.A(_0792_),
    .X(net905));
 sky130_fd_sc_hd__dlygate4sd3_1 hold249 (.A(_0793_),
    .X(net906));
 sky130_fd_sc_hd__dlygate4sd3_1 hold25 (.A(net696),
    .X(net682));
 sky130_fd_sc_hd__dlygate4sd3_1 hold250 (.A(_0380_),
    .X(net907));
 sky130_fd_sc_hd__dlygate4sd3_1 hold251 (.A(la_data_in[26]),
    .X(net908));
 sky130_fd_sc_hd__dlygate4sd3_1 hold252 (.A(net952),
    .X(net909));
 sky130_fd_sc_hd__dlygate4sd3_1 hold253 (.A(net196),
    .X(net910));
 sky130_fd_sc_hd__buf_1 hold254 (.A(_0766_),
    .X(net911));
 sky130_fd_sc_hd__dlygate4sd3_1 hold255 (.A(_0767_),
    .X(net912));
 sky130_fd_sc_hd__dlygate4sd3_1 hold256 (.A(la_data_in[28]),
    .X(net913));
 sky130_fd_sc_hd__dlygate4sd3_1 hold257 (.A(la_data_in[49]),
    .X(net914));
 sky130_fd_sc_hd__dlygate4sd3_1 hold258 (.A(_0403_),
    .X(net915));
 sky130_fd_sc_hd__dlygate4sd3_1 hold259 (.A(net1514),
    .X(net916));
 sky130_fd_sc_hd__buf_8 hold26 (.A(net526),
    .X(net683));
 sky130_fd_sc_hd__dlygate4sd3_1 hold260 (.A(la_data_in[31]),
    .X(net917));
 sky130_fd_sc_hd__dlygate4sd3_1 hold261 (.A(net899),
    .X(net918));
 sky130_fd_sc_hd__dlygate4sd3_1 hold262 (.A(la_data_in[27]),
    .X(net919));
 sky130_fd_sc_hd__dlygate4sd3_1 hold263 (.A(net892),
    .X(net920));
 sky130_fd_sc_hd__dlygate4sd3_1 hold264 (.A(net976),
    .X(net921));
 sky130_fd_sc_hd__dlygate4sd3_1 hold265 (.A(net210),
    .X(net922));
 sky130_fd_sc_hd__buf_1 hold266 (.A(_0742_),
    .X(net923));
 sky130_fd_sc_hd__dlygate4sd3_1 hold267 (.A(_0743_),
    .X(net924));
 sky130_fd_sc_hd__dlygate4sd3_1 hold268 (.A(_0405_),
    .X(net925));
 sky130_fd_sc_hd__dlygate4sd3_1 hold269 (.A(net1081),
    .X(net926));
 sky130_fd_sc_hd__clkbuf_8 hold27 (.A(net521),
    .X(net684));
 sky130_fd_sc_hd__dlygate4sd3_1 hold270 (.A(net242),
    .X(net927));
 sky130_fd_sc_hd__dlygate4sd3_1 hold271 (.A(_0684_),
    .X(net928));
 sky130_fd_sc_hd__dlygate4sd3_1 hold272 (.A(_0685_),
    .X(net929));
 sky130_fd_sc_hd__dlygate4sd3_1 hold273 (.A(_0434_),
    .X(net930));
 sky130_fd_sc_hd__dlygate4sd3_1 hold274 (.A(net935),
    .X(net931));
 sky130_fd_sc_hd__dlygate4sd3_1 hold275 (.A(net187),
    .X(net932));
 sky130_fd_sc_hd__dlymetal6s2s_1 hold276 (.A(_0784_),
    .X(net933));
 sky130_fd_sc_hd__dlygate4sd3_1 hold277 (.A(_0785_),
    .X(net934));
 sky130_fd_sc_hd__dlygate4sd3_1 hold278 (.A(la_data_in[30]),
    .X(net935));
 sky130_fd_sc_hd__dlygate4sd3_1 hold279 (.A(net951),
    .X(net936));
 sky130_fd_sc_hd__dlygate4sd3_1 hold28 (.A(_0356_),
    .X(net685));
 sky130_fd_sc_hd__dlygate4sd3_1 hold280 (.A(net208),
    .X(net937));
 sky130_fd_sc_hd__buf_1 hold281 (.A(_0836_),
    .X(net938));
 sky130_fd_sc_hd__dlygate4sd3_1 hold282 (.A(_0837_),
    .X(net939));
 sky130_fd_sc_hd__dlygate4sd3_1 hold283 (.A(net949),
    .X(net940));
 sky130_fd_sc_hd__dlygate4sd3_1 hold284 (.A(net211),
    .X(net941));
 sky130_fd_sc_hd__buf_1 hold285 (.A(_0740_),
    .X(net942));
 sky130_fd_sc_hd__dlygate4sd3_1 hold286 (.A(_0741_),
    .X(net943));
 sky130_fd_sc_hd__dlygate4sd3_1 hold287 (.A(_0406_),
    .X(net944));
 sky130_fd_sc_hd__dlygate4sd3_1 hold288 (.A(net958),
    .X(net945));
 sky130_fd_sc_hd__dlygate4sd3_1 hold289 (.A(net185),
    .X(net946));
 sky130_fd_sc_hd__dlygate4sd3_1 hold29 (.A(la_data_in[1]),
    .X(net686));
 sky130_fd_sc_hd__dlymetal6s2s_1 hold290 (.A(_0786_),
    .X(net947));
 sky130_fd_sc_hd__dlygate4sd3_1 hold291 (.A(_0912_),
    .X(net948));
 sky130_fd_sc_hd__dlygate4sd3_1 hold292 (.A(la_data_in[52]),
    .X(net949));
 sky130_fd_sc_hd__dlygate4sd3_1 hold293 (.A(_0317_),
    .X(net950));
 sky130_fd_sc_hd__dlygate4sd3_1 hold294 (.A(la_data_in[4]),
    .X(net951));
 sky130_fd_sc_hd__dlygate4sd3_1 hold295 (.A(net1543),
    .X(net952));
 sky130_fd_sc_hd__dlygate4sd3_1 hold296 (.A(net960),
    .X(net953));
 sky130_fd_sc_hd__dlygate4sd3_1 hold297 (.A(net238),
    .X(net954));
 sky130_fd_sc_hd__dlymetal6s2s_1 hold298 (.A(_0690_),
    .X(net955));
 sky130_fd_sc_hd__dlygate4sd3_1 hold299 (.A(_0864_),
    .X(net956));
 sky130_fd_sc_hd__dlygate4sd3_1 hold3 (.A(_0680_),
    .X(net660));
 sky130_fd_sc_hd__dlygate4sd3_1 hold30 (.A(net175),
    .X(net687));
 sky130_fd_sc_hd__dlygate4sd3_1 hold300 (.A(_0342_),
    .X(net957));
 sky130_fd_sc_hd__dlygate4sd3_1 hold301 (.A(net1572),
    .X(net958));
 sky130_fd_sc_hd__dlygate4sd3_1 hold302 (.A(net1559),
    .X(net959));
 sky130_fd_sc_hd__dlygate4sd3_1 hold303 (.A(la_data_in[77]),
    .X(net960));
 sky130_fd_sc_hd__dlygate4sd3_1 hold304 (.A(_0431_),
    .X(net961));
 sky130_fd_sc_hd__dlygate4sd3_1 hold305 (.A(net985),
    .X(net962));
 sky130_fd_sc_hd__dlygate4sd3_1 hold306 (.A(net222),
    .X(net963));
 sky130_fd_sc_hd__buf_1 hold307 (.A(_0720_),
    .X(net964));
 sky130_fd_sc_hd__dlygate4sd3_1 hold308 (.A(_0879_),
    .X(net965));
 sky130_fd_sc_hd__dlygate4sd3_1 hold309 (.A(_0327_),
    .X(net966));
 sky130_fd_sc_hd__dlygate4sd3_1 hold31 (.A(_0842_),
    .X(net688));
 sky130_fd_sc_hd__dlygate4sd3_1 hold310 (.A(net987),
    .X(net967));
 sky130_fd_sc_hd__dlygate4sd3_1 hold311 (.A(net226),
    .X(net968));
 sky130_fd_sc_hd__buf_1 hold312 (.A(_0712_),
    .X(net969));
 sky130_fd_sc_hd__dlygate4sd3_1 hold313 (.A(_0713_),
    .X(net970));
 sky130_fd_sc_hd__dlygate4sd3_1 hold314 (.A(_0420_),
    .X(net971));
 sky130_fd_sc_hd__dlygate4sd3_1 hold315 (.A(net978),
    .X(net972));
 sky130_fd_sc_hd__dlygate4sd3_1 hold316 (.A(net224),
    .X(net973));
 sky130_fd_sc_hd__buf_1 hold317 (.A(_0716_),
    .X(net974));
 sky130_fd_sc_hd__dlygate4sd3_1 hold318 (.A(_0717_),
    .X(net975));
 sky130_fd_sc_hd__dlygate4sd3_1 hold319 (.A(la_data_in[51]),
    .X(net976));
 sky130_fd_sc_hd__dlygate4sd3_1 hold32 (.A(_0940_),
    .X(net689));
 sky130_fd_sc_hd__dlygate4sd3_1 hold320 (.A(_0316_),
    .X(net977));
 sky130_fd_sc_hd__dlygate4sd3_1 hold321 (.A(la_data_in[64]),
    .X(net978));
 sky130_fd_sc_hd__dlygate4sd3_1 hold322 (.A(_0329_),
    .X(net979));
 sky130_fd_sc_hd__dlygate4sd3_1 hold323 (.A(net989),
    .X(net980));
 sky130_fd_sc_hd__dlygate4sd3_1 hold324 (.A(net225),
    .X(net981));
 sky130_fd_sc_hd__buf_1 hold325 (.A(_0714_),
    .X(net982));
 sky130_fd_sc_hd__dlygate4sd3_1 hold326 (.A(_0715_),
    .X(net983));
 sky130_fd_sc_hd__dlygate4sd3_1 hold327 (.A(_0419_),
    .X(net984));
 sky130_fd_sc_hd__dlygate4sd3_1 hold328 (.A(la_data_in[62]),
    .X(net985));
 sky130_fd_sc_hd__dlygate4sd3_1 hold329 (.A(_0416_),
    .X(net986));
 sky130_fd_sc_hd__dlygate4sd3_1 hold33 (.A(_0266_),
    .X(net690));
 sky130_fd_sc_hd__dlygate4sd3_1 hold330 (.A(la_data_in[66]),
    .X(net987));
 sky130_fd_sc_hd__dlygate4sd3_1 hold331 (.A(_0331_),
    .X(net988));
 sky130_fd_sc_hd__dlygate4sd3_1 hold332 (.A(la_data_in[65]),
    .X(net989));
 sky130_fd_sc_hd__dlygate4sd3_1 hold333 (.A(_0330_),
    .X(net990));
 sky130_fd_sc_hd__dlygate4sd3_1 hold334 (.A(net1021),
    .X(net991));
 sky130_fd_sc_hd__dlygate4sd3_1 hold335 (.A(net194),
    .X(net992));
 sky130_fd_sc_hd__buf_1 hold336 (.A(_0770_),
    .X(net993));
 sky130_fd_sc_hd__dlygate4sd3_1 hold337 (.A(_0771_),
    .X(net994));
 sky130_fd_sc_hd__dlygate4sd3_1 hold338 (.A(net1013),
    .X(net995));
 sky130_fd_sc_hd__dlygate4sd3_1 hold339 (.A(net216),
    .X(net996));
 sky130_fd_sc_hd__dlygate4sd3_1 hold34 (.A(la_data_in[82]),
    .X(net691));
 sky130_fd_sc_hd__clkdlybuf4s25_1 hold340 (.A(_0730_),
    .X(net997));
 sky130_fd_sc_hd__dlygate4sd3_1 hold341 (.A(_0731_),
    .X(net998));
 sky130_fd_sc_hd__dlygate4sd3_1 hold342 (.A(net1033),
    .X(net999));
 sky130_fd_sc_hd__dlygate4sd3_1 hold343 (.A(net193),
    .X(net1000));
 sky130_fd_sc_hd__buf_1 hold344 (.A(_0772_),
    .X(net1001));
 sky130_fd_sc_hd__dlygate4sd3_1 hold345 (.A(_0905_),
    .X(net1002));
 sky130_fd_sc_hd__dlygate4sd3_1 hold346 (.A(net1019),
    .X(net1003));
 sky130_fd_sc_hd__dlygate4sd3_1 hold347 (.A(net233),
    .X(net1004));
 sky130_fd_sc_hd__clkbuf_2 hold348 (.A(_0700_),
    .X(net1005));
 sky130_fd_sc_hd__dlygate4sd3_1 hold349 (.A(_0869_),
    .X(net1006));
 sky130_fd_sc_hd__dlymetal6s2s_1 hold35 (.A(net244),
    .X(net692));
 sky130_fd_sc_hd__dlygate4sd3_1 hold350 (.A(_0337_),
    .X(net1007));
 sky130_fd_sc_hd__dlygate4sd3_1 hold351 (.A(net1022),
    .X(net1008));
 sky130_fd_sc_hd__dlygate4sd3_1 hold352 (.A(net212),
    .X(net1009));
 sky130_fd_sc_hd__buf_1 hold353 (.A(_0738_),
    .X(net1010));
 sky130_fd_sc_hd__dlygate4sd3_1 hold354 (.A(_0739_),
    .X(net1011));
 sky130_fd_sc_hd__dlygate4sd3_1 hold355 (.A(_0407_),
    .X(net1012));
 sky130_fd_sc_hd__dlygate4sd3_1 hold356 (.A(la_data_in[57]),
    .X(net1013));
 sky130_fd_sc_hd__dlygate4sd3_1 hold357 (.A(net1044),
    .X(net1014));
 sky130_fd_sc_hd__dlygate4sd3_1 hold358 (.A(net228),
    .X(net1015));
 sky130_fd_sc_hd__buf_1 hold359 (.A(_0708_),
    .X(net1016));
 sky130_fd_sc_hd__dlymetal6s2s_1 hold36 (.A(_0543_),
    .X(net693));
 sky130_fd_sc_hd__dlygate4sd3_1 hold360 (.A(_0709_),
    .X(net1017));
 sky130_fd_sc_hd__dlygate4sd3_1 hold361 (.A(_0422_),
    .X(net1018));
 sky130_fd_sc_hd__dlygate4sd3_1 hold362 (.A(la_data_in[72]),
    .X(net1019));
 sky130_fd_sc_hd__dlygate4sd3_1 hold363 (.A(_0426_),
    .X(net1020));
 sky130_fd_sc_hd__dlygate4sd3_1 hold364 (.A(net1544),
    .X(net1021));
 sky130_fd_sc_hd__dlygate4sd3_1 hold365 (.A(la_data_in[53]),
    .X(net1022));
 sky130_fd_sc_hd__dlygate4sd3_1 hold366 (.A(_0318_),
    .X(net1023));
 sky130_fd_sc_hd__dlygate4sd3_1 hold367 (.A(net1032),
    .X(net1024));
 sky130_fd_sc_hd__dlygate4sd3_1 hold368 (.A(net192),
    .X(net1025));
 sky130_fd_sc_hd__buf_1 hold369 (.A(_0774_),
    .X(net1026));
 sky130_fd_sc_hd__dlygate4sd3_1 hold37 (.A(_0550_),
    .X(net694));
 sky130_fd_sc_hd__dlygate4sd3_1 hold370 (.A(_0906_),
    .X(net1027));
 sky130_fd_sc_hd__dlygate4sd3_1 hold371 (.A(net1154),
    .X(net1028));
 sky130_fd_sc_hd__dlygate4sd3_1 hold372 (.A(net221),
    .X(net1029));
 sky130_fd_sc_hd__dlymetal6s2s_1 hold373 (.A(_0722_),
    .X(net1030));
 sky130_fd_sc_hd__dlygate4sd3_1 hold374 (.A(_0723_),
    .X(net1031));
 sky130_fd_sc_hd__dlygate4sd3_1 hold375 (.A(net1569),
    .X(net1032));
 sky130_fd_sc_hd__dlygate4sd3_1 hold376 (.A(net1565),
    .X(net1033));
 sky130_fd_sc_hd__dlygate4sd3_1 hold377 (.A(net1052),
    .X(net1034));
 sky130_fd_sc_hd__dlygate4sd3_1 hold378 (.A(net227),
    .X(net1035));
 sky130_fd_sc_hd__buf_1 hold379 (.A(_0710_),
    .X(net1036));
 sky130_fd_sc_hd__clkbuf_2 hold38 (.A(net1441),
    .X(net695));
 sky130_fd_sc_hd__dlygate4sd3_1 hold380 (.A(_0874_),
    .X(net1037));
 sky130_fd_sc_hd__dlygate4sd3_1 hold381 (.A(_0332_),
    .X(net1038));
 sky130_fd_sc_hd__dlygate4sd3_1 hold382 (.A(net1054),
    .X(net1039));
 sky130_fd_sc_hd__dlygate4sd3_1 hold383 (.A(net232),
    .X(net1040));
 sky130_fd_sc_hd__buf_1 hold384 (.A(_0702_),
    .X(net1041));
 sky130_fd_sc_hd__dlygate4sd3_1 hold385 (.A(_0870_),
    .X(net1042));
 sky130_fd_sc_hd__dlygate4sd3_1 hold386 (.A(_0336_),
    .X(net1043));
 sky130_fd_sc_hd__dlygate4sd3_1 hold387 (.A(la_data_in[68]),
    .X(net1044));
 sky130_fd_sc_hd__dlygate4sd3_1 hold388 (.A(_0333_),
    .X(net1045));
 sky130_fd_sc_hd__dlygate4sd3_1 hold389 (.A(net1051),
    .X(net1046));
 sky130_fd_sc_hd__dlygate4sd3_1 hold39 (.A(_0683_),
    .X(net696));
 sky130_fd_sc_hd__dlygate4sd3_1 hold390 (.A(net214),
    .X(net1047));
 sky130_fd_sc_hd__buf_1 hold391 (.A(_0734_),
    .X(net1048));
 sky130_fd_sc_hd__dlygate4sd3_1 hold392 (.A(_0886_),
    .X(net1049));
 sky130_fd_sc_hd__dlygate4sd3_1 hold393 (.A(_0320_),
    .X(net1050));
 sky130_fd_sc_hd__dlygate4sd3_1 hold394 (.A(net1540),
    .X(net1051));
 sky130_fd_sc_hd__dlygate4sd3_1 hold395 (.A(la_data_in[67]),
    .X(net1052));
 sky130_fd_sc_hd__dlygate4sd3_1 hold396 (.A(_0421_),
    .X(net1053));
 sky130_fd_sc_hd__dlygate4sd3_1 hold397 (.A(la_data_in[71]),
    .X(net1054));
 sky130_fd_sc_hd__dlygate4sd3_1 hold398 (.A(_0425_),
    .X(net1055));
 sky130_fd_sc_hd__dlygate4sd3_1 hold399 (.A(net1096),
    .X(net1056));
 sky130_fd_sc_hd__dlygate4sd3_1 hold4 (.A(_0435_),
    .X(net661));
 sky130_fd_sc_hd__dlygate4sd3_1 hold40 (.A(net682),
    .X(net697));
 sky130_fd_sc_hd__dlygate4sd3_1 hold400 (.A(net213),
    .X(net1057));
 sky130_fd_sc_hd__buf_1 hold401 (.A(_0736_),
    .X(net1058));
 sky130_fd_sc_hd__dlygate4sd3_1 hold402 (.A(_0887_),
    .X(net1059));
 sky130_fd_sc_hd__dlygate4sd3_1 hold403 (.A(_0319_),
    .X(net1060));
 sky130_fd_sc_hd__dlygate4sd3_1 hold404 (.A(net1113),
    .X(net1061));
 sky130_fd_sc_hd__dlygate4sd3_1 hold405 (.A(net189),
    .X(net1062));
 sky130_fd_sc_hd__dlymetal6s2s_1 hold406 (.A(_0780_),
    .X(net1063));
 sky130_fd_sc_hd__dlygate4sd3_1 hold407 (.A(_0909_),
    .X(net1064));
 sky130_fd_sc_hd__dlygate4sd3_1 hold408 (.A(net1075),
    .X(net1065));
 sky130_fd_sc_hd__dlygate4sd3_1 hold409 (.A(net231),
    .X(net1066));
 sky130_fd_sc_hd__dlygate4sd3_1 hold41 (.A(_0355_),
    .X(net698));
 sky130_fd_sc_hd__buf_1 hold410 (.A(_0704_),
    .X(net1067));
 sky130_fd_sc_hd__dlygate4sd3_1 hold411 (.A(_0871_),
    .X(net1068));
 sky130_fd_sc_hd__dlygate4sd3_1 hold412 (.A(_0335_),
    .X(net1069));
 sky130_fd_sc_hd__dlygate4sd3_1 hold413 (.A(net1137),
    .X(net1070));
 sky130_fd_sc_hd__dlygate4sd3_1 hold414 (.A(net237),
    .X(net1071));
 sky130_fd_sc_hd__dlymetal6s2s_1 hold415 (.A(_0692_),
    .X(net1072));
 sky130_fd_sc_hd__dlygate4sd3_1 hold416 (.A(_0693_),
    .X(net1073));
 sky130_fd_sc_hd__dlygate4sd3_1 hold417 (.A(_0430_),
    .X(net1074));
 sky130_fd_sc_hd__dlygate4sd3_1 hold418 (.A(la_data_in[70]),
    .X(net1075));
 sky130_fd_sc_hd__dlygate4sd3_1 hold419 (.A(_0424_),
    .X(net1076));
 sky130_fd_sc_hd__dlygate4sd3_1 hold42 (.A(net816),
    .X(net699));
 sky130_fd_sc_hd__dlygate4sd3_1 hold420 (.A(net1103),
    .X(net1077));
 sky130_fd_sc_hd__dlygate4sd3_1 hold421 (.A(net234),
    .X(net1078));
 sky130_fd_sc_hd__clkbuf_2 hold422 (.A(_0698_),
    .X(net1079));
 sky130_fd_sc_hd__dlygate4sd3_1 hold423 (.A(_0868_),
    .X(net1080));
 sky130_fd_sc_hd__dlygate4sd3_1 hold424 (.A(la_data_in[80]),
    .X(net1081));
 sky130_fd_sc_hd__dlygate4sd3_1 hold425 (.A(_0345_),
    .X(net1082));
 sky130_fd_sc_hd__dlygate4sd3_1 hold426 (.A(la_data_in[89]),
    .X(net1083));
 sky130_fd_sc_hd__buf_1 hold427 (.A(net251),
    .X(net1084));
 sky130_fd_sc_hd__clkdlybuf4s25_1 hold428 (.A(_0546_),
    .X(net1085));
 sky130_fd_sc_hd__dlygate4sd3_1 hold429 (.A(_0551_),
    .X(net1086));
 sky130_fd_sc_hd__dlygate4sd3_1 hold43 (.A(net201),
    .X(net700));
 sky130_fd_sc_hd__dlygate4sd3_1 hold430 (.A(_0582_),
    .X(net1087));
 sky130_fd_sc_hd__buf_1 hold431 (.A(net1220),
    .X(net1088));
 sky130_fd_sc_hd__dlygate4sd3_1 hold432 (.A(_0856_),
    .X(net1089));
 sky130_fd_sc_hd__dlygate4sd3_1 hold433 (.A(_0349_),
    .X(net1090));
 sky130_fd_sc_hd__dlygate4sd3_1 hold434 (.A(net1111),
    .X(net1091));
 sky130_fd_sc_hd__dlygate4sd3_1 hold435 (.A(net229),
    .X(net1092));
 sky130_fd_sc_hd__buf_1 hold436 (.A(_0706_),
    .X(net1093));
 sky130_fd_sc_hd__dlygate4sd3_1 hold437 (.A(_0872_),
    .X(net1094));
 sky130_fd_sc_hd__dlygate4sd3_1 hold438 (.A(_0334_),
    .X(net1095));
 sky130_fd_sc_hd__dlygate4sd3_1 hold439 (.A(la_data_in[54]),
    .X(net1096));
 sky130_fd_sc_hd__buf_1 hold44 (.A(_0758_),
    .X(net701));
 sky130_fd_sc_hd__dlygate4sd3_1 hold440 (.A(_0408_),
    .X(net1097));
 sky130_fd_sc_hd__dlygate4sd3_1 hold441 (.A(net1116),
    .X(net1098));
 sky130_fd_sc_hd__dlygate4sd3_1 hold442 (.A(net235),
    .X(net1099));
 sky130_fd_sc_hd__dlymetal6s2s_1 hold443 (.A(_0696_),
    .X(net1100));
 sky130_fd_sc_hd__dlygate4sd3_1 hold444 (.A(_0697_),
    .X(net1101));
 sky130_fd_sc_hd__dlygate4sd3_1 hold445 (.A(_0428_),
    .X(net1102));
 sky130_fd_sc_hd__dlygate4sd3_1 hold446 (.A(la_data_in[73]),
    .X(net1103));
 sky130_fd_sc_hd__dlygate4sd3_1 hold447 (.A(_0427_),
    .X(net1104));
 sky130_fd_sc_hd__buf_1 hold448 (.A(net1109),
    .X(net1105));
 sky130_fd_sc_hd__dlygate4sd3_1 hold449 (.A(net215),
    .X(net1106));
 sky130_fd_sc_hd__dlygate4sd3_1 hold45 (.A(_0759_),
    .X(net702));
 sky130_fd_sc_hd__buf_1 hold450 (.A(_0732_),
    .X(net1107));
 sky130_fd_sc_hd__dlygate4sd3_1 hold451 (.A(_0733_),
    .X(net1108));
 sky130_fd_sc_hd__dlygate4sd3_1 hold452 (.A(la_data_in[56]),
    .X(net1109));
 sky130_fd_sc_hd__dlygate4sd3_1 hold453 (.A(_0321_),
    .X(net1110));
 sky130_fd_sc_hd__dlygate4sd3_1 hold454 (.A(la_data_in[69]),
    .X(net1111));
 sky130_fd_sc_hd__dlygate4sd3_1 hold455 (.A(_0423_),
    .X(net1112));
 sky130_fd_sc_hd__dlygate4sd3_1 hold456 (.A(la_data_in[32]),
    .X(net1113));
 sky130_fd_sc_hd__dlygate4sd3_1 hold457 (.A(la_data_in[19]),
    .X(net1114));
 sky130_fd_sc_hd__dlygate4sd3_1 hold458 (.A(net658),
    .X(net1115));
 sky130_fd_sc_hd__dlygate4sd3_1 hold459 (.A(la_data_in[74]),
    .X(net1116));
 sky130_fd_sc_hd__dlygate4sd3_1 hold46 (.A(_0397_),
    .X(net703));
 sky130_fd_sc_hd__dlygate4sd3_1 hold460 (.A(_0339_),
    .X(net1117));
 sky130_fd_sc_hd__dlygate4sd3_1 hold461 (.A(net1123),
    .X(net1118));
 sky130_fd_sc_hd__dlygate4sd3_1 hold462 (.A(net218),
    .X(net1119));
 sky130_fd_sc_hd__dlygate4sd3_1 hold463 (.A(_0726_),
    .X(net1120));
 sky130_fd_sc_hd__dlygate4sd3_1 hold464 (.A(_0882_),
    .X(net1121));
 sky130_fd_sc_hd__dlygate4sd3_1 hold465 (.A(_0324_),
    .X(net1122));
 sky130_fd_sc_hd__dlygate4sd3_1 hold466 (.A(la_data_in[59]),
    .X(net1123));
 sky130_fd_sc_hd__dlygate4sd3_1 hold467 (.A(_0413_),
    .X(net1124));
 sky130_fd_sc_hd__dlygate4sd3_1 hold468 (.A(net1139),
    .X(net1125));
 sky130_fd_sc_hd__dlygate4sd3_1 hold469 (.A(net217),
    .X(net1126));
 sky130_fd_sc_hd__dlygate4sd3_1 hold47 (.A(net807),
    .X(net704));
 sky130_fd_sc_hd__dlygate4sd3_1 hold470 (.A(_0728_),
    .X(net1127));
 sky130_fd_sc_hd__dlygate4sd3_1 hold471 (.A(_0883_),
    .X(net1128));
 sky130_fd_sc_hd__dlygate4sd3_1 hold472 (.A(_0323_),
    .X(net1129));
 sky130_fd_sc_hd__dlygate4sd3_1 hold473 (.A(net1135),
    .X(net1130));
 sky130_fd_sc_hd__dlygate4sd3_1 hold474 (.A(net223),
    .X(net1131));
 sky130_fd_sc_hd__clkdlybuf4s25_1 hold475 (.A(_0718_),
    .X(net1132));
 sky130_fd_sc_hd__dlygate4sd3_1 hold476 (.A(_0878_),
    .X(net1133));
 sky130_fd_sc_hd__dlygate4sd3_1 hold477 (.A(_0328_),
    .X(net1134));
 sky130_fd_sc_hd__dlygate4sd3_1 hold478 (.A(la_data_in[63]),
    .X(net1135));
 sky130_fd_sc_hd__dlygate4sd3_1 hold479 (.A(_0417_),
    .X(net1136));
 sky130_fd_sc_hd__dlygate4sd3_1 hold48 (.A(net164),
    .X(net705));
 sky130_fd_sc_hd__dlygate4sd3_1 hold480 (.A(la_data_in[76]),
    .X(net1137));
 sky130_fd_sc_hd__dlygate4sd3_1 hold481 (.A(_0341_),
    .X(net1138));
 sky130_fd_sc_hd__dlygate4sd3_1 hold482 (.A(la_data_in[58]),
    .X(net1139));
 sky130_fd_sc_hd__dlygate4sd3_1 hold483 (.A(_0412_),
    .X(net1140));
 sky130_fd_sc_hd__dlygate4sd3_1 hold484 (.A(la_data_in[87]),
    .X(net1141));
 sky130_fd_sc_hd__dlygate4sd3_1 hold485 (.A(net249),
    .X(net1142));
 sky130_fd_sc_hd__dlygate4sd3_1 hold486 (.A(_0849_),
    .X(net1143));
 sky130_fd_sc_hd__dlygate4sd3_1 hold487 (.A(_0851_),
    .X(net1144));
 sky130_fd_sc_hd__dlygate4sd3_1 hold488 (.A(_0853_),
    .X(net1145));
 sky130_fd_sc_hd__dlygate4sd3_1 hold489 (.A(_0351_),
    .X(net1146));
 sky130_fd_sc_hd__buf_1 hold49 (.A(_0844_),
    .X(net706));
 sky130_fd_sc_hd__dlygate4sd3_1 hold490 (.A(la_data_in[83]),
    .X(net1147));
 sky130_fd_sc_hd__dlymetal6s2s_1 hold491 (.A(net245),
    .X(net1148));
 sky130_fd_sc_hd__dlygate4sd3_1 hold492 (.A(_0533_),
    .X(net1149));
 sky130_fd_sc_hd__dlygate4sd3_1 hold493 (.A(_0539_),
    .X(net1150));
 sky130_fd_sc_hd__dlygate4sd3_1 hold494 (.A(_0586_),
    .X(net1151));
 sky130_fd_sc_hd__dlygate4sd3_1 hold495 (.A(_0675_),
    .X(net1152));
 sky130_fd_sc_hd__dlygate4sd3_1 hold496 (.A(net1437),
    .X(net1153));
 sky130_fd_sc_hd__dlygate4sd3_1 hold497 (.A(la_data_in[61]),
    .X(net1154));
 sky130_fd_sc_hd__clkdlybuf4s25_1 hold498 (.A(net1162),
    .X(net1155));
 sky130_fd_sc_hd__dlygate4sd3_1 hold499 (.A(net220),
    .X(net1156));
 sky130_fd_sc_hd__dlygate4sd3_1 hold5 (.A(la_data_in[81]),
    .X(net662));
 sky130_fd_sc_hd__dlygate4sd3_1 hold50 (.A(_0941_),
    .X(net707));
 sky130_fd_sc_hd__buf_1 hold500 (.A(_0724_),
    .X(net1157));
 sky130_fd_sc_hd__dlygate4sd3_1 hold501 (.A(_0725_),
    .X(net1158));
 sky130_fd_sc_hd__dlygate4sd3_1 hold502 (.A(_0414_),
    .X(net1159));
 sky130_fd_sc_hd__dlygate4sd3_1 hold503 (.A(la_data_in[18]),
    .X(net1160));
 sky130_fd_sc_hd__dlygate4sd3_1 hold504 (.A(net744),
    .X(net1161));
 sky130_fd_sc_hd__dlygate4sd3_1 hold505 (.A(la_data_in[60]),
    .X(net1162));
 sky130_fd_sc_hd__dlygate4sd3_1 hold506 (.A(_0325_),
    .X(net1163));
 sky130_fd_sc_hd__dlygate4sd3_1 hold507 (.A(la_data_in[17]),
    .X(net1164));
 sky130_fd_sc_hd__dlygate4sd3_1 hold508 (.A(net776),
    .X(net1165));
 sky130_fd_sc_hd__dlygate4sd3_1 hold509 (.A(net1430),
    .X(net1166));
 sky130_fd_sc_hd__dlygate4sd3_1 hold51 (.A(_0265_),
    .X(net708));
 sky130_fd_sc_hd__buf_1 hold510 (.A(net171),
    .X(net1167));
 sky130_fd_sc_hd__dlygate4sd3_1 hold511 (.A(_0521_),
    .X(net1168));
 sky130_fd_sc_hd__buf_1 hold512 (.A(_0812_),
    .X(net1169));
 sky130_fd_sc_hd__dlygate4sd3_1 hold513 (.A(net1174),
    .X(net1170));
 sky130_fd_sc_hd__dlygate4sd3_1 hold514 (.A(net236),
    .X(net1171));
 sky130_fd_sc_hd__dlymetal6s2s_1 hold515 (.A(_0694_),
    .X(net1172));
 sky130_fd_sc_hd__dlygate4sd3_1 hold516 (.A(_0866_),
    .X(net1173));
 sky130_fd_sc_hd__dlygate4sd3_1 hold517 (.A(la_data_in[75]),
    .X(net1174));
 sky130_fd_sc_hd__dlygate4sd3_1 hold518 (.A(_0429_),
    .X(net1175));
 sky130_fd_sc_hd__dlygate4sd3_1 hold519 (.A(net1188),
    .X(net1176));
 sky130_fd_sc_hd__dlygate4sd3_1 hold52 (.A(net830),
    .X(net709));
 sky130_fd_sc_hd__dlygate4sd3_1 hold520 (.A(net176),
    .X(net1177));
 sky130_fd_sc_hd__dlymetal6s2s_1 hold521 (.A(_0804_),
    .X(net1178));
 sky130_fd_sc_hd__dlygate4sd3_1 hold522 (.A(_0805_),
    .X(net1179));
 sky130_fd_sc_hd__dlygate4sd3_1 hold523 (.A(net1190),
    .X(net1180));
 sky130_fd_sc_hd__dlygate4sd3_1 hold524 (.A(net178),
    .X(net1181));
 sky130_fd_sc_hd__dlymetal6s2s_1 hold525 (.A(_0800_),
    .X(net1182));
 sky130_fd_sc_hd__dlygate4sd3_1 hold526 (.A(_0919_),
    .X(net1183));
 sky130_fd_sc_hd__dlygate4sd3_1 hold527 (.A(net1189),
    .X(net1184));
 sky130_fd_sc_hd__dlygate4sd3_1 hold528 (.A(net177),
    .X(net1185));
 sky130_fd_sc_hd__dlymetal6s2s_1 hold529 (.A(_0802_),
    .X(net1186));
 sky130_fd_sc_hd__dlygate4sd3_1 hold53 (.A(net165),
    .X(net710));
 sky130_fd_sc_hd__dlygate4sd3_1 hold530 (.A(_0920_),
    .X(net1187));
 sky130_fd_sc_hd__dlygate4sd3_1 hold531 (.A(la_data_in[20]),
    .X(net1188));
 sky130_fd_sc_hd__dlygate4sd3_1 hold532 (.A(la_data_in[21]),
    .X(net1189));
 sky130_fd_sc_hd__dlygate4sd3_1 hold533 (.A(la_data_in[22]),
    .X(net1190));
 sky130_fd_sc_hd__dlygate4sd3_1 hold534 (.A(net1195),
    .X(net1191));
 sky130_fd_sc_hd__dlygate4sd3_1 hold535 (.A(net179),
    .X(net1192));
 sky130_fd_sc_hd__buf_1 hold536 (.A(_0798_),
    .X(net1193));
 sky130_fd_sc_hd__dlygate4sd3_1 hold537 (.A(_0799_),
    .X(net1194));
 sky130_fd_sc_hd__dlygate4sd3_1 hold538 (.A(la_data_in[23]),
    .X(net1195));
 sky130_fd_sc_hd__dlygate4sd3_1 hold539 (.A(la_data_in[86]),
    .X(net1196));
 sky130_fd_sc_hd__buf_1 hold54 (.A(_0824_),
    .X(net711));
 sky130_fd_sc_hd__dlygate4sd3_1 hold540 (.A(net248),
    .X(net1197));
 sky130_fd_sc_hd__buf_2 hold541 (.A(_0530_),
    .X(net1198));
 sky130_fd_sc_hd__buf_1 hold542 (.A(_0541_),
    .X(net1199));
 sky130_fd_sc_hd__buf_1 hold543 (.A(_0552_),
    .X(net1200));
 sky130_fd_sc_hd__dlygate4sd3_1 hold544 (.A(_0353_),
    .X(net1201));
 sky130_fd_sc_hd__dlygate4sd3_1 hold545 (.A(la_data_in[88]),
    .X(net1202));
 sky130_fd_sc_hd__dlygate4sd3_1 hold546 (.A(net250),
    .X(net1203));
 sky130_fd_sc_hd__dlygate4sd3_1 hold547 (.A(_0547_),
    .X(net1204));
 sky130_fd_sc_hd__dlygate4sd3_1 hold548 (.A(_0548_),
    .X(net1205));
 sky130_fd_sc_hd__dlygate4sd3_1 hold549 (.A(_0562_),
    .X(net1206));
 sky130_fd_sc_hd__dlygate4sd3_1 hold55 (.A(_0931_),
    .X(net712));
 sky130_fd_sc_hd__dlygate4sd3_1 hold550 (.A(net1417),
    .X(net1207));
 sky130_fd_sc_hd__dlygate4sd3_1 hold551 (.A(la_data_in[91]),
    .X(net1208));
 sky130_fd_sc_hd__buf_1 hold552 (.A(net254),
    .X(net1209));
 sky130_fd_sc_hd__dlygate4sd3_1 hold553 (.A(_0558_),
    .X(net1210));
 sky130_fd_sc_hd__dlygate4sd3_1 hold554 (.A(_0559_),
    .X(net1211));
 sky130_fd_sc_hd__dlygate4sd3_1 hold555 (.A(_0676_),
    .X(net1212));
 sky130_fd_sc_hd__dlymetal6s2s_1 hold556 (.A(_0677_),
    .X(net1213));
 sky130_fd_sc_hd__dlygate4sd3_1 hold557 (.A(_0437_),
    .X(net1214));
 sky130_fd_sc_hd__dlygate4sd3_1 hold558 (.A(la_data_in[84]),
    .X(net1215));
 sky130_fd_sc_hd__dlygate4sd3_1 hold559 (.A(net246),
    .X(net1216));
 sky130_fd_sc_hd__dlygate4sd3_1 hold56 (.A(_0275_),
    .X(net713));
 sky130_fd_sc_hd__dlygate4sd3_1 hold560 (.A(_0531_),
    .X(net1217));
 sky130_fd_sc_hd__buf_1 hold561 (.A(_0532_),
    .X(net1218));
 sky130_fd_sc_hd__buf_1 hold562 (.A(net1436),
    .X(net1219));
 sky130_fd_sc_hd__dlygate4sd3_1 hold563 (.A(_0587_),
    .X(net1220));
 sky130_fd_sc_hd__clkbuf_2 hold564 (.A(net1088),
    .X(net1221));
 sky130_fd_sc_hd__dlygate4sd3_1 hold565 (.A(_0461_),
    .X(net1222));
 sky130_fd_sc_hd__dlymetal6s2s_1 hold566 (.A(net1334),
    .X(net1223));
 sky130_fd_sc_hd__clkbuf_2 hold567 (.A(net1335),
    .X(net1224));
 sky130_fd_sc_hd__clkbuf_2 hold568 (.A(net1383),
    .X(net1225));
 sky130_fd_sc_hd__dlygate4sd3_1 hold569 (.A(_0467_),
    .X(net1226));
 sky130_fd_sc_hd__dlygate4sd3_1 hold57 (.A(net856),
    .X(net714));
 sky130_fd_sc_hd__clkbuf_2 hold570 (.A(net1374),
    .X(net1227));
 sky130_fd_sc_hd__dlymetal6s2s_1 hold571 (.A(net1364),
    .X(net1228));
 sky130_fd_sc_hd__clkbuf_2 hold572 (.A(net1346),
    .X(net1229));
 sky130_fd_sc_hd__clkbuf_2 hold573 (.A(net1336),
    .X(net1230));
 sky130_fd_sc_hd__clkbuf_2 hold574 (.A(net1338),
    .X(net1231));
 sky130_fd_sc_hd__dlymetal6s2s_1 hold575 (.A(net1323),
    .X(net1232));
 sky130_fd_sc_hd__clkbuf_2 hold576 (.A(net1361),
    .X(net1233));
 sky130_fd_sc_hd__dlymetal6s2s_1 hold577 (.A(net1371),
    .X(net1234));
 sky130_fd_sc_hd__dlymetal6s2s_1 hold578 (.A(net1321),
    .X(net1235));
 sky130_fd_sc_hd__clkbuf_2 hold579 (.A(net1340),
    .X(net1236));
 sky130_fd_sc_hd__dlygate4sd3_1 hold58 (.A(net204),
    .X(net715));
 sky130_fd_sc_hd__clkbuf_2 hold580 (.A(net1343),
    .X(net1237));
 sky130_fd_sc_hd__buf_1 hold581 (.A(net1378),
    .X(net1238));
 sky130_fd_sc_hd__dlygate4sd3_1 hold582 (.A(_0347_),
    .X(net1239));
 sky130_fd_sc_hd__buf_1 hold583 (.A(net1322),
    .X(net1240));
 sky130_fd_sc_hd__clkbuf_2 hold584 (.A(net1345),
    .X(net1241));
 sky130_fd_sc_hd__dlymetal6s2s_1 hold585 (.A(net1387),
    .X(net1242));
 sky130_fd_sc_hd__clkbuf_2 hold586 (.A(net1358),
    .X(net1243));
 sky130_fd_sc_hd__buf_1 hold587 (.A(net1353),
    .X(net1244));
 sky130_fd_sc_hd__dlymetal6s2s_1 hold588 (.A(net1327),
    .X(net1245));
 sky130_fd_sc_hd__buf_1 hold589 (.A(net1325),
    .X(net1246));
 sky130_fd_sc_hd__dlygate4sd3_1 hold59 (.A(_0752_),
    .X(net716));
 sky130_fd_sc_hd__clkbuf_2 hold590 (.A(net1384),
    .X(net1247));
 sky130_fd_sc_hd__clkbuf_2 hold591 (.A(net1381),
    .X(net1248));
 sky130_fd_sc_hd__dlymetal6s2s_1 hold592 (.A(net1333),
    .X(net1249));
 sky130_fd_sc_hd__dlymetal6s2s_1 hold593 (.A(net1324),
    .X(net1250));
 sky130_fd_sc_hd__buf_1 hold594 (.A(net1355),
    .X(net1251));
 sky130_fd_sc_hd__dlymetal6s2s_1 hold595 (.A(net1331),
    .X(net1252));
 sky130_fd_sc_hd__dlymetal6s2s_1 hold596 (.A(net1342),
    .X(net1253));
 sky130_fd_sc_hd__dlymetal6s2s_1 hold597 (.A(net1376),
    .X(net1254));
 sky130_fd_sc_hd__dlymetal6s2s_1 hold598 (.A(net1365),
    .X(net1255));
 sky130_fd_sc_hd__dlymetal6s2s_1 hold599 (.A(net1389),
    .X(net1256));
 sky130_fd_sc_hd__dlygate4sd3_1 hold6 (.A(net243),
    .X(net663));
 sky130_fd_sc_hd__dlygate4sd3_1 hold60 (.A(_0753_),
    .X(net717));
 sky130_fd_sc_hd__dlymetal6s2s_1 hold600 (.A(net1398),
    .X(net1257));
 sky130_fd_sc_hd__dlygate4sd3_1 hold601 (.A(_0465_),
    .X(net1258));
 sky130_fd_sc_hd__dlymetal6s2s_1 hold602 (.A(net1332),
    .X(net1259));
 sky130_fd_sc_hd__clkbuf_2 hold603 (.A(net1396),
    .X(net1260));
 sky130_fd_sc_hd__clkbuf_2 hold604 (.A(net1392),
    .X(net1261));
 sky130_fd_sc_hd__dlymetal6s2s_1 hold605 (.A(net1385),
    .X(net1262));
 sky130_fd_sc_hd__clkbuf_2 hold606 (.A(net1397),
    .X(net1263));
 sky130_fd_sc_hd__clkbuf_2 hold607 (.A(net1395),
    .X(net1264));
 sky130_fd_sc_hd__buf_1 hold608 (.A(net1393),
    .X(net1265));
 sky130_fd_sc_hd__dlygate4sd3_1 hold609 (.A(_0453_),
    .X(net1266));
 sky130_fd_sc_hd__dlygate4sd3_1 hold61 (.A(_0400_),
    .X(net718));
 sky130_fd_sc_hd__buf_1 hold610 (.A(net1390),
    .X(net1267));
 sky130_fd_sc_hd__dlygate4sd3_1 hold611 (.A(_0463_),
    .X(net1268));
 sky130_fd_sc_hd__buf_1 hold612 (.A(net1388),
    .X(net1269));
 sky130_fd_sc_hd__dlygate4sd3_1 hold613 (.A(_0469_),
    .X(net1270));
 sky130_fd_sc_hd__dlymetal6s2s_1 hold614 (.A(net1382),
    .X(net1271));
 sky130_fd_sc_hd__buf_1 hold615 (.A(net1377),
    .X(net1272));
 sky130_fd_sc_hd__buf_1 hold616 (.A(net1367),
    .X(net1273));
 sky130_fd_sc_hd__dlymetal6s2s_1 hold617 (.A(net1375),
    .X(net1274));
 sky130_fd_sc_hd__dlymetal6s2s_1 hold618 (.A(net1362),
    .X(net1275));
 sky130_fd_sc_hd__dlygate4sd3_1 hold619 (.A(_0483_),
    .X(net1276));
 sky130_fd_sc_hd__dlygate4sd3_1 hold62 (.A(net1576),
    .X(net719));
 sky130_fd_sc_hd__dlymetal6s2s_1 hold620 (.A(net1318),
    .X(net1277));
 sky130_fd_sc_hd__buf_1 hold621 (.A(net1328),
    .X(net1278));
 sky130_fd_sc_hd__dlygate4sd3_1 hold622 (.A(_0479_),
    .X(net1279));
 sky130_fd_sc_hd__dlymetal6s2s_1 hold623 (.A(net1348),
    .X(net1280));
 sky130_fd_sc_hd__dlymetal6s2s_1 hold624 (.A(net1351),
    .X(net1281));
 sky130_fd_sc_hd__clkbuf_2 hold625 (.A(net1369),
    .X(net1282));
 sky130_fd_sc_hd__clkbuf_2 hold626 (.A(net1357),
    .X(net1283));
 sky130_fd_sc_hd__clkbuf_2 hold627 (.A(net1380),
    .X(net1284));
 sky130_fd_sc_hd__clkbuf_2 hold628 (.A(net1386),
    .X(net1285));
 sky130_fd_sc_hd__clkbuf_2 hold629 (.A(net1379),
    .X(net1286));
 sky130_fd_sc_hd__dlygate4sd3_1 hold63 (.A(net230),
    .X(net720));
 sky130_fd_sc_hd__buf_1 hold630 (.A(net1394),
    .X(net1287));
 sky130_fd_sc_hd__dlygate4sd3_1 hold631 (.A(_0493_),
    .X(net1288));
 sky130_fd_sc_hd__dlymetal6s2s_1 hold632 (.A(net1352),
    .X(net1289));
 sky130_fd_sc_hd__buf_1 hold633 (.A(net1391),
    .X(net1290));
 sky130_fd_sc_hd__dlygate4sd3_1 hold634 (.A(_0500_),
    .X(net1291));
 sky130_fd_sc_hd__buf_1 hold635 (.A(net1363),
    .X(net1292));
 sky130_fd_sc_hd__dlymetal6s2s_1 hold636 (.A(net1366),
    .X(net1293));
 sky130_fd_sc_hd__buf_1 hold637 (.A(net1347),
    .X(net1294));
 sky130_fd_sc_hd__clkbuf_2 hold638 (.A(net1344),
    .X(net1295));
 sky130_fd_sc_hd__clkbuf_2 hold639 (.A(net1368),
    .X(net1296));
 sky130_fd_sc_hd__dlymetal6s2s_1 hold64 (.A(_0832_),
    .X(net721));
 sky130_fd_sc_hd__clkbuf_2 hold640 (.A(net1350),
    .X(net1297));
 sky130_fd_sc_hd__clkbuf_2 hold641 (.A(net1339),
    .X(net1298));
 sky130_fd_sc_hd__clkbuf_2 hold642 (.A(net1354),
    .X(net1299));
 sky130_fd_sc_hd__buf_1 hold643 (.A(net1319),
    .X(net1300));
 sky130_fd_sc_hd__clkbuf_2 hold644 (.A(net1341),
    .X(net1301));
 sky130_fd_sc_hd__dlymetal6s2s_1 hold645 (.A(net1326),
    .X(net1302));
 sky130_fd_sc_hd__clkbuf_2 hold646 (.A(net1370),
    .X(net1303));
 sky130_fd_sc_hd__clkbuf_2 hold647 (.A(net1373),
    .X(net1304));
 sky130_fd_sc_hd__buf_1 hold648 (.A(net1317),
    .X(net1305));
 sky130_fd_sc_hd__clkbuf_2 hold649 (.A(net1349),
    .X(net1306));
 sky130_fd_sc_hd__dlygate4sd3_1 hold65 (.A(_0833_),
    .X(net722));
 sky130_fd_sc_hd__clkbuf_2 hold650 (.A(net1356),
    .X(net1307));
 sky130_fd_sc_hd__dlymetal6s2s_1 hold651 (.A(net1320),
    .X(net1308));
 sky130_fd_sc_hd__clkbuf_2 hold652 (.A(net1330),
    .X(net1309));
 sky130_fd_sc_hd__dlymetal6s2s_1 hold653 (.A(net1372),
    .X(net1310));
 sky130_fd_sc_hd__dlygate4sd3_1 hold654 (.A(_0490_),
    .X(net1311));
 sky130_fd_sc_hd__clkbuf_2 hold655 (.A(net1316),
    .X(net1312));
 sky130_fd_sc_hd__buf_1 hold656 (.A(net1337),
    .X(net1313));
 sky130_fd_sc_hd__dlygate4sd3_1 hold657 (.A(_0492_),
    .X(net1314));
 sky130_fd_sc_hd__clkbuf_2 hold658 (.A(net1329),
    .X(net1315));
 sky130_fd_sc_hd__dlygate4sd3_1 hold659 (.A(net1451),
    .X(net1316));
 sky130_fd_sc_hd__dlygate4sd3_1 hold66 (.A(net749),
    .X(net723));
 sky130_fd_sc_hd__dlygate4sd3_1 hold660 (.A(net1459),
    .X(net1317));
 sky130_fd_sc_hd__dlygate4sd3_1 hold661 (.A(net1533),
    .X(net1318));
 sky130_fd_sc_hd__dlygate4sd3_1 hold662 (.A(net1462),
    .X(net1319));
 sky130_fd_sc_hd__dlygate4sd3_1 hold663 (.A(net1505),
    .X(net1320));
 sky130_fd_sc_hd__dlygate4sd3_1 hold664 (.A(net1484),
    .X(net1321));
 sky130_fd_sc_hd__dlygate4sd3_1 hold665 (.A(net1460),
    .X(net1322));
 sky130_fd_sc_hd__dlygate4sd3_1 hold666 (.A(net1485),
    .X(net1323));
 sky130_fd_sc_hd__dlygate4sd3_1 hold667 (.A(net1560),
    .X(net1324));
 sky130_fd_sc_hd__dlygate4sd3_1 hold668 (.A(net1465),
    .X(net1325));
 sky130_fd_sc_hd__dlygate4sd3_1 hold669 (.A(net1520),
    .X(net1326));
 sky130_fd_sc_hd__dlygate4sd3_1 hold67 (.A(net219),
    .X(net724));
 sky130_fd_sc_hd__dlygate4sd3_1 hold670 (.A(net1523),
    .X(net1327));
 sky130_fd_sc_hd__dlygate4sd3_1 hold671 (.A(net1491),
    .X(net1328));
 sky130_fd_sc_hd__dlygate4sd3_1 hold672 (.A(net1468),
    .X(net1329));
 sky130_fd_sc_hd__dlygate4sd3_1 hold673 (.A(net1452),
    .X(net1330));
 sky130_fd_sc_hd__dlygate4sd3_1 hold674 (.A(net1510),
    .X(net1331));
 sky130_fd_sc_hd__dlygate4sd3_1 hold675 (.A(net1508),
    .X(net1332));
 sky130_fd_sc_hd__dlygate4sd3_1 hold676 (.A(net1509),
    .X(net1333));
 sky130_fd_sc_hd__dlygate4sd3_1 hold677 (.A(net1503),
    .X(net1334));
 sky130_fd_sc_hd__dlygate4sd3_1 hold678 (.A(net1457),
    .X(net1335));
 sky130_fd_sc_hd__dlygate4sd3_1 hold679 (.A(net1464),
    .X(net1336));
 sky130_fd_sc_hd__buf_1 hold68 (.A(_0834_),
    .X(net725));
 sky130_fd_sc_hd__dlygate4sd3_1 hold680 (.A(net1480),
    .X(net1337));
 sky130_fd_sc_hd__dlygate4sd3_1 hold681 (.A(net1469),
    .X(net1338));
 sky130_fd_sc_hd__dlygate4sd3_1 hold682 (.A(net1455),
    .X(net1339));
 sky130_fd_sc_hd__dlygate4sd3_1 hold683 (.A(net1458),
    .X(net1340));
 sky130_fd_sc_hd__dlygate4sd3_1 hold684 (.A(net1467),
    .X(net1341));
 sky130_fd_sc_hd__dlygate4sd3_1 hold685 (.A(net1506),
    .X(net1342));
 sky130_fd_sc_hd__dlygate4sd3_1 hold686 (.A(net1466),
    .X(net1343));
 sky130_fd_sc_hd__dlygate4sd3_1 hold687 (.A(net1456),
    .X(net1344));
 sky130_fd_sc_hd__dlygate4sd3_1 hold688 (.A(net1453),
    .X(net1345));
 sky130_fd_sc_hd__dlygate4sd3_1 hold689 (.A(net1471),
    .X(net1346));
 sky130_fd_sc_hd__dlygate4sd3_1 hold69 (.A(_0835_),
    .X(net726));
 sky130_fd_sc_hd__dlygate4sd3_1 hold690 (.A(net1482),
    .X(net1347));
 sky130_fd_sc_hd__dlygate4sd3_1 hold691 (.A(net1519),
    .X(net1348));
 sky130_fd_sc_hd__dlygate4sd3_1 hold692 (.A(net1479),
    .X(net1349));
 sky130_fd_sc_hd__dlygate4sd3_1 hold693 (.A(net1470),
    .X(net1350));
 sky130_fd_sc_hd__dlygate4sd3_1 hold694 (.A(net1521),
    .X(net1351));
 sky130_fd_sc_hd__dlygate4sd3_1 hold695 (.A(net1564),
    .X(net1352));
 sky130_fd_sc_hd__dlygate4sd3_1 hold696 (.A(net1486),
    .X(net1353));
 sky130_fd_sc_hd__dlygate4sd3_1 hold697 (.A(net1477),
    .X(net1354));
 sky130_fd_sc_hd__dlygate4sd3_1 hold698 (.A(net1504),
    .X(net1355));
 sky130_fd_sc_hd__dlygate4sd3_1 hold699 (.A(net1472),
    .X(net1356));
 sky130_fd_sc_hd__dlygate4sd3_1 hold7 (.A(_0859_),
    .X(net664));
 sky130_fd_sc_hd__dlygate4sd3_1 hold70 (.A(net837),
    .X(net727));
 sky130_fd_sc_hd__dlygate4sd3_1 hold700 (.A(net1463),
    .X(net1357));
 sky130_fd_sc_hd__dlygate4sd3_1 hold701 (.A(net1494),
    .X(net1358));
 sky130_fd_sc_hd__dlygate4sd3_1 hold702 (.A(net1419),
    .X(net1359));
 sky130_fd_sc_hd__buf_12 hold703 (.A(net1360),
    .X(la_data_out[113]));
 sky130_fd_sc_hd__dlygate4sd3_1 hold704 (.A(net1474),
    .X(net1361));
 sky130_fd_sc_hd__dlygate4sd3_1 hold705 (.A(net1550),
    .X(net1362));
 sky130_fd_sc_hd__dlygate4sd3_1 hold706 (.A(net1511),
    .X(net1363));
 sky130_fd_sc_hd__dlygate4sd3_1 hold707 (.A(net1553),
    .X(net1364));
 sky130_fd_sc_hd__dlygate4sd3_1 hold708 (.A(net1522),
    .X(net1365));
 sky130_fd_sc_hd__dlygate4sd3_1 hold709 (.A(net1562),
    .X(net1366));
 sky130_fd_sc_hd__dlygate4sd3_1 hold71 (.A(net200),
    .X(net728));
 sky130_fd_sc_hd__dlygate4sd3_1 hold710 (.A(net1493),
    .X(net1367));
 sky130_fd_sc_hd__dlygate4sd3_1 hold711 (.A(net1476),
    .X(net1368));
 sky130_fd_sc_hd__dlygate4sd3_1 hold712 (.A(net1483),
    .X(net1369));
 sky130_fd_sc_hd__dlygate4sd3_1 hold713 (.A(net1478),
    .X(net1370));
 sky130_fd_sc_hd__dlygate4sd3_1 hold714 (.A(net1563),
    .X(net1371));
 sky130_fd_sc_hd__dlygate4sd3_1 hold715 (.A(net1528),
    .X(net1372));
 sky130_fd_sc_hd__dlygate4sd3_1 hold716 (.A(net1488),
    .X(net1373));
 sky130_fd_sc_hd__dlygate4sd3_1 hold717 (.A(net1475),
    .X(net1374));
 sky130_fd_sc_hd__dlygate4sd3_1 hold718 (.A(net1529),
    .X(net1375));
 sky130_fd_sc_hd__dlygate4sd3_1 hold719 (.A(net1537),
    .X(net1376));
 sky130_fd_sc_hd__buf_1 hold72 (.A(_0760_),
    .X(net729));
 sky130_fd_sc_hd__dlygate4sd3_1 hold720 (.A(net1513),
    .X(net1377));
 sky130_fd_sc_hd__dlygate4sd3_1 hold721 (.A(net1517),
    .X(net1378));
 sky130_fd_sc_hd__dlygate4sd3_1 hold722 (.A(net1481),
    .X(net1379));
 sky130_fd_sc_hd__dlygate4sd3_1 hold723 (.A(net1487),
    .X(net1380));
 sky130_fd_sc_hd__dlygate4sd3_1 hold724 (.A(net1490),
    .X(net1381));
 sky130_fd_sc_hd__dlygate4sd3_1 hold725 (.A(net1534),
    .X(net1382));
 sky130_fd_sc_hd__dlygate4sd3_1 hold726 (.A(net1512),
    .X(net1383));
 sky130_fd_sc_hd__dlygate4sd3_1 hold727 (.A(net1502),
    .X(net1384));
 sky130_fd_sc_hd__dlygate4sd3_1 hold728 (.A(net1524),
    .X(net1385));
 sky130_fd_sc_hd__dlygate4sd3_1 hold729 (.A(net1473),
    .X(net1386));
 sky130_fd_sc_hd__dlygate4sd3_1 hold73 (.A(_0761_),
    .X(net730));
 sky130_fd_sc_hd__dlygate4sd3_1 hold730 (.A(net1554),
    .X(net1387));
 sky130_fd_sc_hd__dlygate4sd3_1 hold731 (.A(net1507),
    .X(net1388));
 sky130_fd_sc_hd__dlygate4sd3_1 hold732 (.A(net1542),
    .X(net1389));
 sky130_fd_sc_hd__dlygate4sd3_1 hold733 (.A(net1516),
    .X(net1390));
 sky130_fd_sc_hd__dlygate4sd3_1 hold734 (.A(net1525),
    .X(net1391));
 sky130_fd_sc_hd__dlygate4sd3_1 hold735 (.A(net1495),
    .X(net1392));
 sky130_fd_sc_hd__dlygate4sd3_1 hold736 (.A(net1518),
    .X(net1393));
 sky130_fd_sc_hd__dlygate4sd3_1 hold737 (.A(net1532),
    .X(net1394));
 sky130_fd_sc_hd__dlygate4sd3_1 hold738 (.A(net1489),
    .X(net1395));
 sky130_fd_sc_hd__dlygate4sd3_1 hold739 (.A(net1492),
    .X(net1396));
 sky130_fd_sc_hd__dlygate4sd3_1 hold74 (.A(_0396_),
    .X(net731));
 sky130_fd_sc_hd__dlygate4sd3_1 hold740 (.A(net1496),
    .X(net1397));
 sky130_fd_sc_hd__dlygate4sd3_1 hold741 (.A(net1568),
    .X(net1398));
 sky130_fd_sc_hd__dlygate4sd3_1 hold742 (.A(net1421),
    .X(net1399));
 sky130_fd_sc_hd__buf_12 hold743 (.A(net1400),
    .X(la_data_out[54]));
 sky130_fd_sc_hd__buf_1 hold744 (.A(net1422),
    .X(net1401));
 sky130_fd_sc_hd__buf_12 hold745 (.A(net1402),
    .X(la_data_out[123]));
 sky130_fd_sc_hd__dlygate4sd3_1 hold746 (.A(net1420),
    .X(net1403));
 sky130_fd_sc_hd__buf_12 hold747 (.A(net1404),
    .X(la_data_out[73]));
 sky130_fd_sc_hd__buf_1 hold748 (.A(net1424),
    .X(net1405));
 sky130_fd_sc_hd__buf_12 hold749 (.A(net1406),
    .X(la_data_out[122]));
 sky130_fd_sc_hd__dlygate4sd3_1 hold75 (.A(la_data_in[93]),
    .X(net732));
 sky130_fd_sc_hd__buf_1 hold750 (.A(net1426),
    .X(net1407));
 sky130_fd_sc_hd__buf_12 hold751 (.A(net1408),
    .X(la_data_out[125]));
 sky130_fd_sc_hd__buf_1 hold752 (.A(net1428),
    .X(net1409));
 sky130_fd_sc_hd__buf_12 hold753 (.A(net1410),
    .X(la_data_out[124]));
 sky130_fd_sc_hd__dlygate4sd3_1 hold754 (.A(net1434),
    .X(net1411));
 sky130_fd_sc_hd__dlygate4sd3_1 hold755 (.A(_0534_),
    .X(net1412));
 sky130_fd_sc_hd__dlygate4sd3_1 hold756 (.A(_0848_),
    .X(net1413));
 sky130_fd_sc_hd__dlygate4sd3_1 hold757 (.A(_0352_),
    .X(net1414));
 sky130_fd_sc_hd__dlygate4sd3_1 hold758 (.A(net1442),
    .X(net1415));
 sky130_fd_sc_hd__dlygate4sd3_1 hold759 (.A(_0561_),
    .X(net1416));
 sky130_fd_sc_hd__dlymetal6s2s_1 hold76 (.A(net256),
    .X(net733));
 sky130_fd_sc_hd__dlygate4sd3_1 hold760 (.A(_0436_),
    .X(net1417));
 sky130_fd_sc_hd__dlygate4sd3_1 hold761 (.A(net1438),
    .X(net1418));
 sky130_fd_sc_hd__dlygate4sd3_1 hold762 (.A(net440),
    .X(net1419));
 sky130_fd_sc_hd__dlygate4sd3_1 hold763 (.A(net488),
    .X(net1420));
 sky130_fd_sc_hd__dlygate4sd3_1 hold764 (.A(net469),
    .X(net1421));
 sky130_fd_sc_hd__dlygate4sd3_1 hold765 (.A(net442),
    .X(net1422));
 sky130_fd_sc_hd__dlygate4sd3_1 hold766 (.A(net1401),
    .X(net1423));
 sky130_fd_sc_hd__dlygate4sd3_1 hold767 (.A(net441),
    .X(net1424));
 sky130_fd_sc_hd__dlygate4sd3_1 hold768 (.A(net1405),
    .X(net1425));
 sky130_fd_sc_hd__dlygate4sd3_1 hold769 (.A(net444),
    .X(net1426));
 sky130_fd_sc_hd__dlygate4sd3_1 hold77 (.A(_0580_),
    .X(net734));
 sky130_fd_sc_hd__dlygate4sd3_1 hold770 (.A(net1407),
    .X(net1427));
 sky130_fd_sc_hd__dlygate4sd3_1 hold771 (.A(net443),
    .X(net1428));
 sky130_fd_sc_hd__dlygate4sd3_1 hold772 (.A(net1409),
    .X(net1429));
 sky130_fd_sc_hd__dlygate4sd3_1 hold773 (.A(la_data_in[16]),
    .X(net1430));
 sky130_fd_sc_hd__dlygate4sd3_1 hold774 (.A(_0281_),
    .X(net1431));
 sky130_fd_sc_hd__dlygate4sd3_1 hold775 (.A(\reg_temp[98] ),
    .X(net1432));
 sky130_fd_sc_hd__dlygate4sd3_1 hold776 (.A(\reg_temp[75] ),
    .X(net1433));
 sky130_fd_sc_hd__dlygate4sd3_1 hold777 (.A(la_data_in[85]),
    .X(net1434));
 sky130_fd_sc_hd__dlygate4sd3_1 hold778 (.A(_0584_),
    .X(net1435));
 sky130_fd_sc_hd__dlygate4sd3_1 hold779 (.A(_0585_),
    .X(net1436));
 sky130_fd_sc_hd__dlygate4sd3_1 hold78 (.A(_0581_),
    .X(net735));
 sky130_fd_sc_hd__dlygate4sd3_1 hold780 (.A(_0438_),
    .X(net1437));
 sky130_fd_sc_hd__dlygate4sd3_1 hold781 (.A(la_data_in[90]),
    .X(net1438));
 sky130_fd_sc_hd__dlygate4sd3_1 hold782 (.A(_0555_),
    .X(net1439));
 sky130_fd_sc_hd__dlygate4sd3_1 hold783 (.A(_0556_),
    .X(net1440));
 sky130_fd_sc_hd__dlygate4sd3_1 hold784 (.A(_0560_),
    .X(net1441));
 sky130_fd_sc_hd__dlygate4sd3_1 hold785 (.A(la_data_in[92]),
    .X(net1442));
 sky130_fd_sc_hd__dlygate4sd3_1 hold786 (.A(\reg_temp[39] ),
    .X(net1443));
 sky130_fd_sc_hd__dlygate4sd3_1 hold787 (.A(\reg_temp[131] ),
    .X(net1444));
 sky130_fd_sc_hd__dlygate4sd3_1 hold788 (.A(\reg_temp[79] ),
    .X(net1445));
 sky130_fd_sc_hd__dlygate4sd3_1 hold789 (.A(_0595_),
    .X(net1446));
 sky130_fd_sc_hd__clkbuf_2 hold79 (.A(net769),
    .X(net736));
 sky130_fd_sc_hd__dlygate4sd3_1 hold790 (.A(\reg_temp[80] ),
    .X(net1447));
 sky130_fd_sc_hd__dlygate4sd3_1 hold791 (.A(_0594_),
    .X(net1448));
 sky130_fd_sc_hd__dlygate4sd3_1 hold792 (.A(\reg_temp[46] ),
    .X(net1449));
 sky130_fd_sc_hd__dlygate4sd3_1 hold793 (.A(\reg_temp[38] ),
    .X(net1450));
 sky130_fd_sc_hd__dlygate4sd3_1 hold794 (.A(net448),
    .X(net1451));
 sky130_fd_sc_hd__dlygate4sd3_1 hold795 (.A(net499),
    .X(net1452));
 sky130_fd_sc_hd__dlygate4sd3_1 hold796 (.A(net485),
    .X(net1453));
 sky130_fd_sc_hd__dlygate4sd3_1 hold797 (.A(\reg_temp[43] ),
    .X(net1454));
 sky130_fd_sc_hd__dlygate4sd3_1 hold798 (.A(net459),
    .X(net1455));
 sky130_fd_sc_hd__dlygate4sd3_1 hold799 (.A(net455),
    .X(net1456));
 sky130_fd_sc_hd__dlygate4sd3_1 hold8 (.A(_0860_),
    .X(net665));
 sky130_fd_sc_hd__buf_6 hold80 (.A(net537),
    .X(net737));
 sky130_fd_sc_hd__dlygate4sd3_1 hold800 (.A(net463),
    .X(net1457));
 sky130_fd_sc_hd__dlygate4sd3_1 hold801 (.A(net495),
    .X(net1458));
 sky130_fd_sc_hd__dlygate4sd3_1 hold802 (.A(net482),
    .X(net1459));
 sky130_fd_sc_hd__dlygate4sd3_1 hold803 (.A(net439),
    .X(net1460));
 sky130_fd_sc_hd__dlygate4sd3_1 hold804 (.A(la_data_in[2]),
    .X(net1461));
 sky130_fd_sc_hd__dlygate4sd3_1 hold805 (.A(net481),
    .X(net1462));
 sky130_fd_sc_hd__dlygate4sd3_1 hold806 (.A(net466),
    .X(net1463));
 sky130_fd_sc_hd__dlygate4sd3_1 hold807 (.A(net512),
    .X(net1464));
 sky130_fd_sc_hd__dlygate4sd3_1 hold808 (.A(net513),
    .X(net1465));
 sky130_fd_sc_hd__dlygate4sd3_1 hold809 (.A(net497),
    .X(net1466));
 sky130_fd_sc_hd__buf_4 hold81 (.A(net536),
    .X(net738));
 sky130_fd_sc_hd__dlygate4sd3_1 hold810 (.A(net511),
    .X(net1467));
 sky130_fd_sc_hd__dlygate4sd3_1 hold811 (.A(net453),
    .X(net1468));
 sky130_fd_sc_hd__dlygate4sd3_1 hold812 (.A(net496),
    .X(net1469));
 sky130_fd_sc_hd__dlygate4sd3_1 hold813 (.A(net460),
    .X(net1470));
 sky130_fd_sc_hd__dlygate4sd3_1 hold814 (.A(net493),
    .X(net1471));
 sky130_fd_sc_hd__dlygate4sd3_1 hold815 (.A(net431),
    .X(net1472));
 sky130_fd_sc_hd__dlygate4sd3_1 hold816 (.A(net451),
    .X(net1473));
 sky130_fd_sc_hd__dlygate4sd3_1 hold817 (.A(net507),
    .X(net1474));
 sky130_fd_sc_hd__dlygate4sd3_1 hold818 (.A(net465),
    .X(net1475));
 sky130_fd_sc_hd__dlygate4sd3_1 hold819 (.A(net467),
    .X(net1476));
 sky130_fd_sc_hd__dlygate4sd3_1 hold82 (.A(_0271_),
    .X(net739));
 sky130_fd_sc_hd__dlygate4sd3_1 hold820 (.A(net479),
    .X(net1477));
 sky130_fd_sc_hd__dlygate4sd3_1 hold821 (.A(net484),
    .X(net1478));
 sky130_fd_sc_hd__dlygate4sd3_1 hold822 (.A(net483),
    .X(net1479));
 sky130_fd_sc_hd__dlygate4sd3_1 hold823 (.A(net500),
    .X(net1480));
 sky130_fd_sc_hd__dlygate4sd3_1 hold824 (.A(net458),
    .X(net1481));
 sky130_fd_sc_hd__dlygate4sd3_1 hold825 (.A(net435),
    .X(net1482));
 sky130_fd_sc_hd__dlygate4sd3_1 hold826 (.A(net450),
    .X(net1483));
 sky130_fd_sc_hd__dlygate4sd3_1 hold827 (.A(net510),
    .X(net1484));
 sky130_fd_sc_hd__dlygate4sd3_1 hold828 (.A(net506),
    .X(net1485));
 sky130_fd_sc_hd__dlygate4sd3_1 hold829 (.A(net437),
    .X(net1486));
 sky130_fd_sc_hd__dlygate4sd3_1 hold83 (.A(net755),
    .X(net740));
 sky130_fd_sc_hd__dlygate4sd3_1 hold830 (.A(net457),
    .X(net1487));
 sky130_fd_sc_hd__dlygate4sd3_1 hold831 (.A(net480),
    .X(net1488));
 sky130_fd_sc_hd__dlygate4sd3_1 hold832 (.A(net464),
    .X(net1489));
 sky130_fd_sc_hd__dlygate4sd3_1 hold833 (.A(net427),
    .X(net1490));
 sky130_fd_sc_hd__dlygate4sd3_1 hold834 (.A(net487),
    .X(net1491));
 sky130_fd_sc_hd__dlygate4sd3_1 hold835 (.A(net449),
    .X(net1492));
 sky130_fd_sc_hd__dlygate4sd3_1 hold836 (.A(net470),
    .X(net1493));
 sky130_fd_sc_hd__dlygate4sd3_1 hold837 (.A(net494),
    .X(net1494));
 sky130_fd_sc_hd__dlygate4sd3_1 hold838 (.A(net452),
    .X(net1495));
 sky130_fd_sc_hd__dlygate4sd3_1 hold839 (.A(net462),
    .X(net1496));
 sky130_fd_sc_hd__dlygate4sd3_1 hold84 (.A(net169),
    .X(net741));
 sky130_fd_sc_hd__dlygate4sd3_1 hold840 (.A(la_data_in[0]),
    .X(net1497));
 sky130_fd_sc_hd__dlygate4sd3_1 hold841 (.A(_0354_),
    .X(net1498));
 sky130_fd_sc_hd__dlygate4sd3_1 hold842 (.A(la_data_in[12]),
    .X(net1499));
 sky130_fd_sc_hd__dlygate4sd3_1 hold843 (.A(_0366_),
    .X(net1500));
 sky130_fd_sc_hd__dlygate4sd3_1 hold844 (.A(la_data_in[43]),
    .X(net1501));
 sky130_fd_sc_hd__dlygate4sd3_1 hold845 (.A(net514),
    .X(net1502));
 sky130_fd_sc_hd__dlygate4sd3_1 hold846 (.A(net492),
    .X(net1503));
 sky130_fd_sc_hd__dlygate4sd3_1 hold847 (.A(net429),
    .X(net1504));
 sky130_fd_sc_hd__dlygate4sd3_1 hold848 (.A(net509),
    .X(net1505));
 sky130_fd_sc_hd__dlygate4sd3_1 hold849 (.A(net432),
    .X(net1506));
 sky130_fd_sc_hd__buf_1 hold85 (.A(_0816_),
    .X(net742));
 sky130_fd_sc_hd__dlygate4sd3_1 hold850 (.A(net477),
    .X(net1507));
 sky130_fd_sc_hd__dlygate4sd3_1 hold851 (.A(net433),
    .X(net1508));
 sky130_fd_sc_hd__dlygate4sd3_1 hold852 (.A(net428),
    .X(net1509));
 sky130_fd_sc_hd__dlygate4sd3_1 hold853 (.A(net430),
    .X(net1510));
 sky130_fd_sc_hd__dlygate4sd3_1 hold854 (.A(net502),
    .X(net1511));
 sky130_fd_sc_hd__dlygate4sd3_1 hold855 (.A(net475),
    .X(net1512));
 sky130_fd_sc_hd__dlygate4sd3_1 hold856 (.A(net478),
    .X(net1513));
 sky130_fd_sc_hd__dlygate4sd3_1 hold857 (.A(la_data_in[44]),
    .X(net1514));
 sky130_fd_sc_hd__dlygate4sd3_1 hold858 (.A(_0309_),
    .X(net1515));
 sky130_fd_sc_hd__dlygate4sd3_1 hold859 (.A(net471),
    .X(net1516));
 sky130_fd_sc_hd__dlygate4sd3_1 hold86 (.A(_0817_),
    .X(net743));
 sky130_fd_sc_hd__dlygate4sd3_1 hold860 (.A(net445),
    .X(net1517));
 sky130_fd_sc_hd__dlygate4sd3_1 hold861 (.A(net461),
    .X(net1518));
 sky130_fd_sc_hd__dlygate4sd3_1 hold862 (.A(net454),
    .X(net1519));
 sky130_fd_sc_hd__dlygate4sd3_1 hold863 (.A(net505),
    .X(net1520));
 sky130_fd_sc_hd__dlygate4sd3_1 hold864 (.A(net456),
    .X(net1521));
 sky130_fd_sc_hd__dlygate4sd3_1 hold865 (.A(net476),
    .X(net1522));
 sky130_fd_sc_hd__dlygate4sd3_1 hold866 (.A(net438),
    .X(net1523));
 sky130_fd_sc_hd__dlygate4sd3_1 hold867 (.A(net447),
    .X(net1524));
 sky130_fd_sc_hd__dlygate4sd3_1 hold868 (.A(net508),
    .X(net1525));
 sky130_fd_sc_hd__dlygate4sd3_1 hold869 (.A(la_data_in[40]),
    .X(net1526));
 sky130_fd_sc_hd__dlygate4sd3_1 hold87 (.A(net1160),
    .X(net744));
 sky130_fd_sc_hd__dlygate4sd3_1 hold870 (.A(_0394_),
    .X(net1527));
 sky130_fd_sc_hd__dlygate4sd3_1 hold871 (.A(net498),
    .X(net1528));
 sky130_fd_sc_hd__dlygate4sd3_1 hold872 (.A(net468),
    .X(net1529));
 sky130_fd_sc_hd__dlygate4sd3_1 hold873 (.A(la_data_in[9]),
    .X(net1530));
 sky130_fd_sc_hd__dlygate4sd3_1 hold874 (.A(_0363_),
    .X(net1531));
 sky130_fd_sc_hd__dlygate4sd3_1 hold875 (.A(net501),
    .X(net1532));
 sky130_fd_sc_hd__dlygate4sd3_1 hold876 (.A(net489),
    .X(net1533));
 sky130_fd_sc_hd__dlygate4sd3_1 hold877 (.A(net474),
    .X(net1534));
 sky130_fd_sc_hd__dlygate4sd3_1 hold878 (.A(la_data_in[11]),
    .X(net1535));
 sky130_fd_sc_hd__dlygate4sd3_1 hold879 (.A(_0365_),
    .X(net1536));
 sky130_fd_sc_hd__clkbuf_2 hold88 (.A(net173),
    .X(net745));
 sky130_fd_sc_hd__dlygate4sd3_1 hold880 (.A(net472),
    .X(net1537));
 sky130_fd_sc_hd__dlygate4sd3_1 hold881 (.A(la_data_in[42]),
    .X(net1538));
 sky130_fd_sc_hd__dlygate4sd3_1 hold882 (.A(_0307_),
    .X(net1539));
 sky130_fd_sc_hd__dlygate4sd3_1 hold883 (.A(la_data_in[55]),
    .X(net1540));
 sky130_fd_sc_hd__dlygate4sd3_1 hold884 (.A(_0409_),
    .X(net1541));
 sky130_fd_sc_hd__dlygate4sd3_1 hold885 (.A(net436),
    .X(net1542));
 sky130_fd_sc_hd__dlygate4sd3_1 hold886 (.A(la_data_in[39]),
    .X(net1543));
 sky130_fd_sc_hd__dlygate4sd3_1 hold887 (.A(la_data_in[37]),
    .X(net1544));
 sky130_fd_sc_hd__dlygate4sd3_1 hold888 (.A(_0302_),
    .X(net1545));
 sky130_fd_sc_hd__dlygate4sd3_1 hold889 (.A(la_data_in[14]),
    .X(net1546));
 sky130_fd_sc_hd__dlygate4sd3_1 hold89 (.A(_0847_),
    .X(net746));
 sky130_fd_sc_hd__dlygate4sd3_1 hold890 (.A(_0279_),
    .X(net1547));
 sky130_fd_sc_hd__dlygate4sd3_1 hold891 (.A(la_data_in[41]),
    .X(net1548));
 sky130_fd_sc_hd__dlygate4sd3_1 hold892 (.A(_0395_),
    .X(net1549));
 sky130_fd_sc_hd__dlygate4sd3_1 hold893 (.A(net491),
    .X(net1550));
 sky130_fd_sc_hd__dlygate4sd3_1 hold894 (.A(la_data_in[8]),
    .X(net1551));
 sky130_fd_sc_hd__dlygate4sd3_1 hold895 (.A(_0362_),
    .X(net1552));
 sky130_fd_sc_hd__dlygate4sd3_1 hold896 (.A(net434),
    .X(net1553));
 sky130_fd_sc_hd__dlygate4sd3_1 hold897 (.A(net486),
    .X(net1554));
 sky130_fd_sc_hd__dlygate4sd3_1 hold898 (.A(la_data_in[3]),
    .X(net1555));
 sky130_fd_sc_hd__dlygate4sd3_1 hold899 (.A(_0357_),
    .X(net1556));
 sky130_fd_sc_hd__dlygate4sd3_1 hold9 (.A(_0346_),
    .X(net666));
 sky130_fd_sc_hd__dlygate4sd3_1 hold90 (.A(net1413),
    .X(net747));
 sky130_fd_sc_hd__dlygate4sd3_1 hold900 (.A(la_data_in[10]),
    .X(net1557));
 sky130_fd_sc_hd__dlygate4sd3_1 hold901 (.A(_0364_),
    .X(net1558));
 sky130_fd_sc_hd__dlygate4sd3_1 hold902 (.A(la_data_in[38]),
    .X(net1559));
 sky130_fd_sc_hd__dlygate4sd3_1 hold903 (.A(net490),
    .X(net1560));
 sky130_fd_sc_hd__dlygate4sd3_1 hold904 (.A(\reg_temp[146] ),
    .X(net1561));
 sky130_fd_sc_hd__dlygate4sd3_1 hold905 (.A(net504),
    .X(net1562));
 sky130_fd_sc_hd__dlygate4sd3_1 hold906 (.A(net446),
    .X(net1563));
 sky130_fd_sc_hd__dlygate4sd3_1 hold907 (.A(net503),
    .X(net1564));
 sky130_fd_sc_hd__dlygate4sd3_1 hold908 (.A(la_data_in[36]),
    .X(net1565));
 sky130_fd_sc_hd__dlygate4sd3_1 hold909 (.A(_0390_),
    .X(net1566));
 sky130_fd_sc_hd__dlygate4sd3_1 hold91 (.A(net1414),
    .X(net748));
 sky130_fd_sc_hd__dlygate4sd3_1 hold910 (.A(\reg_temp[73] ),
    .X(net1567));
 sky130_fd_sc_hd__dlygate4sd3_1 hold911 (.A(net473),
    .X(net1568));
 sky130_fd_sc_hd__dlygate4sd3_1 hold912 (.A(la_data_in[35]),
    .X(net1569));
 sky130_fd_sc_hd__dlygate4sd3_1 hold913 (.A(_0389_),
    .X(net1570));
 sky130_fd_sc_hd__dlygate4sd3_1 hold914 (.A(\reg_temp[61] ),
    .X(net1571));
 sky130_fd_sc_hd__dlygate4sd3_1 hold915 (.A(la_data_in[29]),
    .X(net1572));
 sky130_fd_sc_hd__dlygate4sd3_1 hold916 (.A(_0383_),
    .X(net1573));
 sky130_fd_sc_hd__dlygate4sd3_1 hold917 (.A(la_data_in[7]),
    .X(net1574));
 sky130_fd_sc_hd__dlygate4sd3_1 hold918 (.A(_0272_),
    .X(net1575));
 sky130_fd_sc_hd__dlygate4sd3_1 hold919 (.A(la_data_in[6]),
    .X(net1576));
 sky130_fd_sc_hd__dlygate4sd3_1 hold92 (.A(la_data_in[5]),
    .X(net749));
 sky130_fd_sc_hd__dlygate4sd3_1 hold920 (.A(_0360_),
    .X(net1577));
 sky130_fd_sc_hd__dlygate4sd3_1 hold921 (.A(\reg_temp[32] ),
    .X(net1578));
 sky130_fd_sc_hd__dlygate4sd3_1 hold922 (.A(\reg_temp[99] ),
    .X(net1579));
 sky130_fd_sc_hd__dlygate4sd3_1 hold923 (.A(\reg_temp[97] ),
    .X(net1580));
 sky130_fd_sc_hd__dlygate4sd3_1 hold924 (.A(\reg_temp[143] ),
    .X(net1581));
 sky130_fd_sc_hd__dlygate4sd3_1 hold925 (.A(\reg_temp[104] ),
    .X(net1582));
 sky130_fd_sc_hd__dlygate4sd3_1 hold926 (.A(\reg_temp[109] ),
    .X(net1583));
 sky130_fd_sc_hd__dlygate4sd3_1 hold927 (.A(\reg_temp[24] ),
    .X(net1584));
 sky130_fd_sc_hd__dlygate4sd3_1 hold928 (.A(_0289_),
    .X(net1585));
 sky130_fd_sc_hd__dlygate4sd3_1 hold929 (.A(\reg_temp[30] ),
    .X(net1586));
 sky130_fd_sc_hd__dlygate4sd3_1 hold93 (.A(net817),
    .X(net750));
 sky130_fd_sc_hd__dlygate4sd3_1 hold930 (.A(\reg_temp[49] ),
    .X(net1587));
 sky130_fd_sc_hd__dlygate4sd3_1 hold931 (.A(\reg_temp[126] ),
    .X(net1588));
 sky130_fd_sc_hd__dlygate4sd3_1 hold932 (.A(\reg_temp[12] ),
    .X(net1589));
 sky130_fd_sc_hd__dlygate4sd3_1 hold933 (.A(\reg_temp[33] ),
    .X(net1590));
 sky130_fd_sc_hd__dlygate4sd3_1 hold934 (.A(_0298_),
    .X(net1591));
 sky130_fd_sc_hd__dlygate4sd3_1 hold935 (.A(\reg_temp[116] ),
    .X(net1592));
 sky130_fd_sc_hd__dlygate4sd3_1 hold936 (.A(_0388_),
    .X(net1593));
 sky130_fd_sc_hd__dlygate4sd3_1 hold937 (.A(\reg_temp[31] ),
    .X(net1594));
 sky130_fd_sc_hd__dlygate4sd3_1 hold938 (.A(\reg_temp[26] ),
    .X(net1595));
 sky130_fd_sc_hd__dlygate4sd3_1 hold939 (.A(_0291_),
    .X(net1596));
 sky130_fd_sc_hd__dlygate4sd3_1 hold94 (.A(net205),
    .X(net751));
 sky130_fd_sc_hd__dlygate4sd3_1 hold940 (.A(\reg_temp[34] ),
    .X(net1597));
 sky130_fd_sc_hd__dlygate4sd3_1 hold941 (.A(\reg_temp[113] ),
    .X(net1598));
 sky130_fd_sc_hd__dlygate4sd3_1 hold942 (.A(\reg_temp[15] ),
    .X(net1599));
 sky130_fd_sc_hd__dlygate4sd3_1 hold943 (.A(_0280_),
    .X(net1600));
 sky130_fd_sc_hd__dlygate4sd3_1 hold944 (.A(\reg_temp[112] ),
    .X(net1601));
 sky130_fd_sc_hd__dlygate4sd3_1 hold945 (.A(\reg_temp[57] ),
    .X(net1602));
 sky130_fd_sc_hd__dlygate4sd3_1 hold946 (.A(_0322_),
    .X(net1603));
 sky130_fd_sc_hd__dlygate4sd3_1 hold947 (.A(\reg_temp[110] ),
    .X(net1604));
 sky130_fd_sc_hd__dlygate4sd3_1 hold948 (.A(\reg_temp[120] ),
    .X(net1605));
 sky130_fd_sc_hd__dlygate4sd3_1 hold949 (.A(\reg_temp[96] ),
    .X(net1606));
 sky130_fd_sc_hd__buf_1 hold95 (.A(_0750_),
    .X(net752));
 sky130_fd_sc_hd__dlygate4sd3_1 hold950 (.A(\reg_temp[36] ),
    .X(net1607));
 sky130_fd_sc_hd__dlygate4sd3_1 hold951 (.A(\reg_temp[4] ),
    .X(net1608));
 sky130_fd_sc_hd__dlygate4sd3_1 hold952 (.A(_0269_),
    .X(net1609));
 sky130_fd_sc_hd__dlygate4sd3_1 hold953 (.A(\reg_temp[95] ),
    .X(net1610));
 sky130_fd_sc_hd__dlygate4sd3_1 hold954 (.A(_0367_),
    .X(net1611));
 sky130_fd_sc_hd__dlygate4sd3_1 hold955 (.A(\reg_temp[103] ),
    .X(net1612));
 sky130_fd_sc_hd__dlygate4sd3_1 hold956 (.A(\reg_temp[27] ),
    .X(net1613));
 sky130_fd_sc_hd__dlygate4sd3_1 hold957 (.A(\reg_temp[138] ),
    .X(net1614));
 sky130_fd_sc_hd__dlygate4sd3_1 hold958 (.A(\reg_temp[5] ),
    .X(net1615));
 sky130_fd_sc_hd__dlygate4sd3_1 hold959 (.A(\reg_temp[114] ),
    .X(net1616));
 sky130_fd_sc_hd__dlygate4sd3_1 hold96 (.A(_0751_),
    .X(net753));
 sky130_fd_sc_hd__dlygate4sd3_1 hold960 (.A(_0386_),
    .X(net1617));
 sky130_fd_sc_hd__dlygate4sd3_1 hold961 (.A(\reg_temp[121] ),
    .X(net1618));
 sky130_fd_sc_hd__dlygate4sd3_1 hold962 (.A(\reg_temp[28] ),
    .X(net1619));
 sky130_fd_sc_hd__dlygate4sd3_1 hold963 (.A(\reg_temp[18] ),
    .X(net1620));
 sky130_fd_sc_hd__dlygate4sd3_1 hold964 (.A(\reg_temp[19] ),
    .X(net1621));
 sky130_fd_sc_hd__dlygate4sd3_1 hold965 (.A(\reg_temp[3] ),
    .X(net1622));
 sky130_fd_sc_hd__dlygate4sd3_1 hold966 (.A(\reg_temp[101] ),
    .X(net1623));
 sky130_fd_sc_hd__dlygate4sd3_1 hold967 (.A(\reg_temp[87] ),
    .X(net1624));
 sky130_fd_sc_hd__dlygate4sd3_1 hold968 (.A(\reg_temp[119] ),
    .X(net1625));
 sky130_fd_sc_hd__dlygate4sd3_1 hold969 (.A(\reg_temp[25] ),
    .X(net1626));
 sky130_fd_sc_hd__dlygate4sd3_1 hold97 (.A(_0401_),
    .X(net754));
 sky130_fd_sc_hd__dlygate4sd3_1 hold970 (.A(\reg_temp[100] ),
    .X(net1627));
 sky130_fd_sc_hd__dlygate4sd3_1 hold971 (.A(\reg_temp[82] ),
    .X(net1628));
 sky130_fd_sc_hd__dlygate4sd3_1 hold972 (.A(\reg_temp[13] ),
    .X(net1629));
 sky130_fd_sc_hd__dlygate4sd3_1 hold973 (.A(\reg_temp[21] ),
    .X(net1630));
 sky130_fd_sc_hd__dlygate4sd3_1 hold974 (.A(\reg_temp[139] ),
    .X(net1631));
 sky130_fd_sc_hd__dlygate4sd3_1 hold975 (.A(\reg_temp[102] ),
    .X(net1632));
 sky130_fd_sc_hd__dlygate4sd3_1 hold976 (.A(\reg_temp[123] ),
    .X(net1633));
 sky130_fd_sc_hd__dlygate4sd3_1 hold977 (.A(\reg_temp[89] ),
    .X(net1634));
 sky130_fd_sc_hd__dlygate4sd3_1 hold978 (.A(\reg_temp[115] ),
    .X(net1635));
 sky130_fd_sc_hd__dlygate4sd3_1 hold979 (.A(\reg_temp[86] ),
    .X(net1636));
 sky130_fd_sc_hd__dlygate4sd3_1 hold98 (.A(net1546),
    .X(net755));
 sky130_fd_sc_hd__dlygate4sd3_1 hold980 (.A(\reg_temp[20] ),
    .X(net1637));
 sky130_fd_sc_hd__dlygate4sd3_1 hold981 (.A(\reg_temp[22] ),
    .X(net1638));
 sky130_fd_sc_hd__dlygate4sd3_1 hold982 (.A(\reg_temp[29] ),
    .X(net1639));
 sky130_fd_sc_hd__dlygate4sd3_1 hold983 (.A(\reg_temp[4] ),
    .X(net1640));
 sky130_fd_sc_hd__dlygate4sd3_1 hold984 (.A(\reg_temp[85] ),
    .X(net1641));
 sky130_fd_sc_hd__dlygate4sd3_1 hold985 (.A(\reg_temp[17] ),
    .X(net1642));
 sky130_fd_sc_hd__dlygate4sd3_1 hold986 (.A(\reg_temp[105] ),
    .X(net1643));
 sky130_fd_sc_hd__dlygate4sd3_1 hold987 (.A(\reg_temp[35] ),
    .X(net1644));
 sky130_fd_sc_hd__dlygate4sd3_1 hold988 (.A(\reg_temp[92] ),
    .X(net1645));
 sky130_fd_sc_hd__dlygate4sd3_1 hold989 (.A(\reg_temp[41] ),
    .X(net1646));
 sky130_fd_sc_hd__dlygate4sd3_1 hold99 (.A(net829),
    .X(net756));
 sky130_fd_sc_hd__dlygate4sd3_1 hold990 (.A(\reg_temp[23] ),
    .X(net1647));
 sky130_fd_sc_hd__dlygate4sd3_1 hold991 (.A(\reg_temp[40] ),
    .X(net1648));
 sky130_fd_sc_hd__dlygate4sd3_1 hold992 (.A(\reg_temp[93] ),
    .X(net1649));
 sky130_fd_sc_hd__dlygate4sd3_1 hold993 (.A(\reg_temp[8] ),
    .X(net1650));
 sky130_fd_sc_hd__dlygate4sd3_1 hold994 (.A(\reg_temp[58] ),
    .X(net1651));
 sky130_fd_sc_hd__buf_1 input1 (.A(data_in[0]),
    .X(net1));
 sky130_fd_sc_hd__clkbuf_1 input10 (.A(data_in[108]),
    .X(net10));
 sky130_fd_sc_hd__buf_1 input100 (.A(data_in[42]),
    .X(net100));
 sky130_fd_sc_hd__buf_1 input101 (.A(data_in[43]),
    .X(net101));
 sky130_fd_sc_hd__buf_1 input102 (.A(data_in[44]),
    .X(net102));
 sky130_fd_sc_hd__buf_1 input103 (.A(data_in[45]),
    .X(net103));
 sky130_fd_sc_hd__dlymetal6s2s_1 input104 (.A(data_in[46]),
    .X(net104));
 sky130_fd_sc_hd__buf_1 input105 (.A(data_in[47]),
    .X(net105));
 sky130_fd_sc_hd__buf_1 input106 (.A(data_in[48]),
    .X(net106));
 sky130_fd_sc_hd__buf_1 input107 (.A(data_in[49]),
    .X(net107));
 sky130_fd_sc_hd__buf_1 input108 (.A(data_in[4]),
    .X(net108));
 sky130_fd_sc_hd__buf_1 input109 (.A(data_in[50]),
    .X(net109));
 sky130_fd_sc_hd__clkbuf_1 input11 (.A(data_in[109]),
    .X(net11));
 sky130_fd_sc_hd__buf_1 input110 (.A(data_in[51]),
    .X(net110));
 sky130_fd_sc_hd__buf_1 input111 (.A(data_in[52]),
    .X(net111));
 sky130_fd_sc_hd__buf_1 input112 (.A(data_in[53]),
    .X(net112));
 sky130_fd_sc_hd__buf_1 input113 (.A(data_in[54]),
    .X(net113));
 sky130_fd_sc_hd__buf_1 input114 (.A(data_in[55]),
    .X(net114));
 sky130_fd_sc_hd__buf_1 input115 (.A(data_in[56]),
    .X(net115));
 sky130_fd_sc_hd__buf_1 input116 (.A(data_in[57]),
    .X(net116));
 sky130_fd_sc_hd__dlymetal6s2s_1 input117 (.A(data_in[58]),
    .X(net117));
 sky130_fd_sc_hd__buf_1 input118 (.A(data_in[59]),
    .X(net118));
 sky130_fd_sc_hd__clkbuf_1 input119 (.A(data_in[5]),
    .X(net119));
 sky130_fd_sc_hd__buf_1 input12 (.A(data_in[10]),
    .X(net12));
 sky130_fd_sc_hd__dlymetal6s2s_1 input120 (.A(data_in[60]),
    .X(net120));
 sky130_fd_sc_hd__clkbuf_2 input121 (.A(data_in[61]),
    .X(net121));
 sky130_fd_sc_hd__clkbuf_2 input122 (.A(data_in[62]),
    .X(net122));
 sky130_fd_sc_hd__clkbuf_2 input123 (.A(data_in[63]),
    .X(net123));
 sky130_fd_sc_hd__clkbuf_2 input124 (.A(data_in[64]),
    .X(net124));
 sky130_fd_sc_hd__clkbuf_2 input125 (.A(data_in[65]),
    .X(net125));
 sky130_fd_sc_hd__clkbuf_2 input126 (.A(data_in[66]),
    .X(net126));
 sky130_fd_sc_hd__buf_2 input127 (.A(data_in[67]),
    .X(net127));
 sky130_fd_sc_hd__buf_2 input128 (.A(data_in[68]),
    .X(net128));
 sky130_fd_sc_hd__clkbuf_2 input129 (.A(data_in[69]),
    .X(net129));
 sky130_fd_sc_hd__clkbuf_1 input13 (.A(data_in[110]),
    .X(net13));
 sky130_fd_sc_hd__clkbuf_1 input130 (.A(data_in[6]),
    .X(net130));
 sky130_fd_sc_hd__clkbuf_2 input131 (.A(data_in[70]),
    .X(net131));
 sky130_fd_sc_hd__clkbuf_2 input132 (.A(data_in[71]),
    .X(net132));
 sky130_fd_sc_hd__clkbuf_2 input133 (.A(data_in[72]),
    .X(net133));
 sky130_fd_sc_hd__buf_2 input134 (.A(data_in[73]),
    .X(net134));
 sky130_fd_sc_hd__buf_2 input135 (.A(data_in[74]),
    .X(net135));
 sky130_fd_sc_hd__clkbuf_2 input136 (.A(data_in[75]),
    .X(net136));
 sky130_fd_sc_hd__clkbuf_2 input137 (.A(data_in[76]),
    .X(net137));
 sky130_fd_sc_hd__buf_2 input138 (.A(data_in[77]),
    .X(net138));
 sky130_fd_sc_hd__buf_2 input139 (.A(data_in[78]),
    .X(net139));
 sky130_fd_sc_hd__clkbuf_1 input14 (.A(data_in[111]),
    .X(net14));
 sky130_fd_sc_hd__buf_2 input140 (.A(data_in[79]),
    .X(net140));
 sky130_fd_sc_hd__clkbuf_1 input141 (.A(data_in[7]),
    .X(net141));
 sky130_fd_sc_hd__dlymetal6s2s_1 input142 (.A(data_in[80]),
    .X(net142));
 sky130_fd_sc_hd__buf_1 input143 (.A(data_in[81]),
    .X(net143));
 sky130_fd_sc_hd__buf_1 input144 (.A(data_in[82]),
    .X(net144));
 sky130_fd_sc_hd__buf_1 input145 (.A(data_in[83]),
    .X(net145));
 sky130_fd_sc_hd__buf_1 input146 (.A(data_in[84]),
    .X(net146));
 sky130_fd_sc_hd__buf_1 input147 (.A(data_in[85]),
    .X(net147));
 sky130_fd_sc_hd__buf_1 input148 (.A(data_in[86]),
    .X(net148));
 sky130_fd_sc_hd__buf_1 input149 (.A(data_in[87]),
    .X(net149));
 sky130_fd_sc_hd__clkbuf_1 input15 (.A(data_in[112]),
    .X(net15));
 sky130_fd_sc_hd__buf_1 input150 (.A(data_in[88]),
    .X(net150));
 sky130_fd_sc_hd__clkbuf_1 input151 (.A(data_in[89]),
    .X(net151));
 sky130_fd_sc_hd__buf_1 input152 (.A(data_in[8]),
    .X(net152));
 sky130_fd_sc_hd__buf_1 input153 (.A(data_in[90]),
    .X(net153));
 sky130_fd_sc_hd__buf_1 input154 (.A(data_in[91]),
    .X(net154));
 sky130_fd_sc_hd__buf_1 input155 (.A(data_in[92]),
    .X(net155));
 sky130_fd_sc_hd__buf_1 input156 (.A(data_in[93]),
    .X(net156));
 sky130_fd_sc_hd__buf_1 input157 (.A(data_in[94]),
    .X(net157));
 sky130_fd_sc_hd__buf_1 input158 (.A(data_in[95]),
    .X(net158));
 sky130_fd_sc_hd__buf_1 input159 (.A(data_in[96]),
    .X(net159));
 sky130_fd_sc_hd__clkbuf_1 input16 (.A(data_in[113]),
    .X(net16));
 sky130_fd_sc_hd__buf_1 input160 (.A(data_in[97]),
    .X(net160));
 sky130_fd_sc_hd__buf_1 input161 (.A(data_in[98]),
    .X(net161));
 sky130_fd_sc_hd__clkbuf_1 input162 (.A(data_in[99]),
    .X(net162));
 sky130_fd_sc_hd__buf_1 input163 (.A(data_in[9]),
    .X(net163));
 sky130_fd_sc_hd__clkbuf_1 input164 (.A(net704),
    .X(net164));
 sky130_fd_sc_hd__clkbuf_1 input165 (.A(net709),
    .X(net165));
 sky130_fd_sc_hd__clkbuf_1 input166 (.A(net811),
    .X(net166));
 sky130_fd_sc_hd__clkbuf_1 input167 (.A(net858),
    .X(net167));
 sky130_fd_sc_hd__buf_1 input168 (.A(net874),
    .X(net168));
 sky130_fd_sc_hd__clkbuf_1 input169 (.A(net740),
    .X(net169));
 sky130_fd_sc_hd__clkbuf_1 input17 (.A(data_in[114]),
    .X(net17));
 sky130_fd_sc_hd__clkbuf_1 input170 (.A(net787),
    .X(net170));
 sky130_fd_sc_hd__buf_1 input171 (.A(net1166),
    .X(net171));
 sky130_fd_sc_hd__buf_1 input172 (.A(net1165),
    .X(net172));
 sky130_fd_sc_hd__buf_1 input173 (.A(net1161),
    .X(net173));
 sky130_fd_sc_hd__buf_1 input174 (.A(net1115),
    .X(net174));
 sky130_fd_sc_hd__clkbuf_1 input175 (.A(net686),
    .X(net175));
 sky130_fd_sc_hd__dlymetal6s2s_1 input176 (.A(net1176),
    .X(net176));
 sky130_fd_sc_hd__dlymetal6s2s_1 input177 (.A(net1184),
    .X(net177));
 sky130_fd_sc_hd__dlymetal6s2s_1 input178 (.A(net1180),
    .X(net178));
 sky130_fd_sc_hd__dlymetal6s2s_1 input179 (.A(net1191),
    .X(net179));
 sky130_fd_sc_hd__clkbuf_1 input18 (.A(data_in[115]),
    .X(net18));
 sky130_fd_sc_hd__clkbuf_1 input180 (.A(net782),
    .X(net180));
 sky130_fd_sc_hd__buf_1 input181 (.A(net863),
    .X(net181));
 sky130_fd_sc_hd__clkbuf_1 input182 (.A(net903),
    .X(net182));
 sky130_fd_sc_hd__clkbuf_1 input183 (.A(net920),
    .X(net183));
 sky130_fd_sc_hd__clkbuf_1 input184 (.A(net878),
    .X(net184));
 sky130_fd_sc_hd__clkbuf_1 input185 (.A(net945),
    .X(net185));
 sky130_fd_sc_hd__clkbuf_1 input186 (.A(net672),
    .X(net186));
 sky130_fd_sc_hd__buf_1 input187 (.A(net931),
    .X(net187));
 sky130_fd_sc_hd__clkbuf_1 input188 (.A(net918),
    .X(net188));
 sky130_fd_sc_hd__buf_1 input189 (.A(net1061),
    .X(net189));
 sky130_fd_sc_hd__clkbuf_1 input19 (.A(data_in[116]),
    .X(net19));
 sky130_fd_sc_hd__clkbuf_1 input190 (.A(net761),
    .X(net190));
 sky130_fd_sc_hd__buf_1 input191 (.A(net791),
    .X(net191));
 sky130_fd_sc_hd__clkbuf_1 input192 (.A(net1024),
    .X(net192));
 sky130_fd_sc_hd__clkbuf_1 input193 (.A(net999),
    .X(net193));
 sky130_fd_sc_hd__clkbuf_1 input194 (.A(net991),
    .X(net194));
 sky130_fd_sc_hd__clkbuf_1 input195 (.A(net882),
    .X(net195));
 sky130_fd_sc_hd__clkbuf_1 input196 (.A(net909),
    .X(net196));
 sky130_fd_sc_hd__clkbuf_1 input197 (.A(net831),
    .X(net197));
 sky130_fd_sc_hd__clkbuf_1 input198 (.A(net846),
    .X(net198));
 sky130_fd_sc_hd__clkbuf_1 input199 (.A(net838),
    .X(net199));
 sky130_fd_sc_hd__clkbuf_1 input2 (.A(data_in[100]),
    .X(net2));
 sky130_fd_sc_hd__clkbuf_1 input20 (.A(data_in[117]),
    .X(net20));
 sky130_fd_sc_hd__clkbuf_1 input200 (.A(net727),
    .X(net200));
 sky130_fd_sc_hd__clkbuf_1 input201 (.A(net699),
    .X(net201));
 sky130_fd_sc_hd__clkbuf_1 input202 (.A(net852),
    .X(net202));
 sky130_fd_sc_hd__clkbuf_1 input203 (.A(net667),
    .X(net203));
 sky130_fd_sc_hd__clkbuf_1 input204 (.A(net714),
    .X(net204));
 sky130_fd_sc_hd__clkbuf_1 input205 (.A(net750),
    .X(net205));
 sky130_fd_sc_hd__clkbuf_1 input206 (.A(net796),
    .X(net206));
 sky130_fd_sc_hd__buf_1 input207 (.A(net802),
    .X(net207));
 sky130_fd_sc_hd__clkbuf_1 input208 (.A(net936),
    .X(net208));
 sky130_fd_sc_hd__clkbuf_1 input209 (.A(net819),
    .X(net209));
 sky130_fd_sc_hd__buf_1 input21 (.A(data_in[118]),
    .X(net21));
 sky130_fd_sc_hd__buf_1 input210 (.A(net921),
    .X(net210));
 sky130_fd_sc_hd__clkbuf_1 input211 (.A(net940),
    .X(net211));
 sky130_fd_sc_hd__buf_1 input212 (.A(net1008),
    .X(net212));
 sky130_fd_sc_hd__clkbuf_1 input213 (.A(net1056),
    .X(net213));
 sky130_fd_sc_hd__clkbuf_1 input214 (.A(net1046),
    .X(net214));
 sky130_fd_sc_hd__clkbuf_1 input215 (.A(net1105),
    .X(net215));
 sky130_fd_sc_hd__buf_1 input216 (.A(net995),
    .X(net216));
 sky130_fd_sc_hd__buf_1 input217 (.A(net1125),
    .X(net217));
 sky130_fd_sc_hd__clkbuf_1 input218 (.A(net1118),
    .X(net218));
 sky130_fd_sc_hd__buf_1 input219 (.A(net723),
    .X(net219));
 sky130_fd_sc_hd__buf_1 input22 (.A(data_in[119]),
    .X(net22));
 sky130_fd_sc_hd__buf_1 input220 (.A(net1155),
    .X(net220));
 sky130_fd_sc_hd__clkbuf_1 input221 (.A(net1028),
    .X(net221));
 sky130_fd_sc_hd__clkbuf_1 input222 (.A(net962),
    .X(net222));
 sky130_fd_sc_hd__buf_1 input223 (.A(net1130),
    .X(net223));
 sky130_fd_sc_hd__clkbuf_1 input224 (.A(net972),
    .X(net224));
 sky130_fd_sc_hd__clkbuf_1 input225 (.A(net980),
    .X(net225));
 sky130_fd_sc_hd__clkbuf_1 input226 (.A(net967),
    .X(net226));
 sky130_fd_sc_hd__clkbuf_1 input227 (.A(net1034),
    .X(net227));
 sky130_fd_sc_hd__clkbuf_1 input228 (.A(net1014),
    .X(net228));
 sky130_fd_sc_hd__clkbuf_1 input229 (.A(net1091),
    .X(net229));
 sky130_fd_sc_hd__buf_1 input23 (.A(data_in[11]),
    .X(net23));
 sky130_fd_sc_hd__buf_1 input230 (.A(net719),
    .X(net230));
 sky130_fd_sc_hd__clkbuf_1 input231 (.A(net1065),
    .X(net231));
 sky130_fd_sc_hd__clkbuf_1 input232 (.A(net1039),
    .X(net232));
 sky130_fd_sc_hd__buf_1 input233 (.A(net1003),
    .X(net233));
 sky130_fd_sc_hd__clkbuf_1 input234 (.A(net1077),
    .X(net234));
 sky130_fd_sc_hd__clkbuf_1 input235 (.A(net1098),
    .X(net235));
 sky130_fd_sc_hd__clkbuf_1 input236 (.A(net1170),
    .X(net236));
 sky130_fd_sc_hd__clkbuf_1 input237 (.A(net1070),
    .X(net237));
 sky130_fd_sc_hd__clkbuf_1 input238 (.A(net953),
    .X(net238));
 sky130_fd_sc_hd__clkbuf_1 input239 (.A(net886),
    .X(net239));
 sky130_fd_sc_hd__buf_1 input24 (.A(data_in[120]),
    .X(net24));
 sky130_fd_sc_hd__clkbuf_1 input240 (.A(net824),
    .X(net240));
 sky130_fd_sc_hd__clkbuf_1 input241 (.A(net772),
    .X(net241));
 sky130_fd_sc_hd__clkbuf_1 input242 (.A(net926),
    .X(net242));
 sky130_fd_sc_hd__clkbuf_1 input243 (.A(net662),
    .X(net243));
 sky130_fd_sc_hd__clkbuf_1 input244 (.A(net691),
    .X(net244));
 sky130_fd_sc_hd__clkbuf_1 input245 (.A(net1147),
    .X(net245));
 sky130_fd_sc_hd__dlymetal6s2s_1 input246 (.A(net1215),
    .X(net246));
 sky130_fd_sc_hd__clkbuf_2 input247 (.A(net1411),
    .X(net247));
 sky130_fd_sc_hd__buf_1 input248 (.A(net1196),
    .X(net248));
 sky130_fd_sc_hd__buf_1 input249 (.A(net1141),
    .X(net249));
 sky130_fd_sc_hd__buf_1 input25 (.A(data_in[121]),
    .X(net25));
 sky130_fd_sc_hd__buf_1 input250 (.A(net1202),
    .X(net250));
 sky130_fd_sc_hd__clkbuf_1 input251 (.A(net1083),
    .X(net251));
 sky130_fd_sc_hd__buf_1 input252 (.A(net842),
    .X(net252));
 sky130_fd_sc_hd__buf_1 input253 (.A(net1418),
    .X(net253));
 sky130_fd_sc_hd__clkbuf_1 input254 (.A(net1208),
    .X(net254));
 sky130_fd_sc_hd__dlymetal6s2s_1 input255 (.A(net1415),
    .X(net255));
 sky130_fd_sc_hd__clkbuf_1 input256 (.A(net732),
    .X(net256));
 sky130_fd_sc_hd__clkbuf_1 input257 (.A(net765),
    .X(net257));
 sky130_fd_sc_hd__clkbuf_1 input258 (.A(net677),
    .X(net258));
 sky130_fd_sc_hd__clkbuf_1 input259 (.A(net756),
    .X(net259));
 sky130_fd_sc_hd__buf_1 input26 (.A(data_in[122]),
    .X(net26));
 sky130_fd_sc_hd__clkbuf_2 input260 (.A(next_key),
    .X(net260));
 sky130_fd_sc_hd__buf_2 input261 (.A(slv_done),
    .X(net261));
 sky130_fd_sc_hd__clkbuf_8 input262 (.A(wb_rst_i),
    .X(net262));
 sky130_fd_sc_hd__buf_1 input27 (.A(data_in[123]),
    .X(net27));
 sky130_fd_sc_hd__buf_1 input28 (.A(data_in[124]),
    .X(net28));
 sky130_fd_sc_hd__buf_1 input29 (.A(data_in[125]),
    .X(net29));
 sky130_fd_sc_hd__clkbuf_1 input3 (.A(data_in[101]),
    .X(net3));
 sky130_fd_sc_hd__buf_1 input30 (.A(data_in[126]),
    .X(net30));
 sky130_fd_sc_hd__buf_1 input31 (.A(data_in[127]),
    .X(net31));
 sky130_fd_sc_hd__buf_1 input32 (.A(data_in[128]),
    .X(net32));
 sky130_fd_sc_hd__buf_1 input33 (.A(data_in[129]),
    .X(net33));
 sky130_fd_sc_hd__buf_1 input34 (.A(data_in[12]),
    .X(net34));
 sky130_fd_sc_hd__buf_1 input35 (.A(data_in[130]),
    .X(net35));
 sky130_fd_sc_hd__buf_1 input36 (.A(data_in[131]),
    .X(net36));
 sky130_fd_sc_hd__buf_1 input37 (.A(data_in[132]),
    .X(net37));
 sky130_fd_sc_hd__buf_1 input38 (.A(data_in[133]),
    .X(net38));
 sky130_fd_sc_hd__buf_1 input39 (.A(data_in[134]),
    .X(net39));
 sky130_fd_sc_hd__clkbuf_1 input4 (.A(data_in[102]),
    .X(net4));
 sky130_fd_sc_hd__clkbuf_1 input40 (.A(data_in[135]),
    .X(net40));
 sky130_fd_sc_hd__clkbuf_1 input41 (.A(data_in[136]),
    .X(net41));
 sky130_fd_sc_hd__clkbuf_1 input42 (.A(data_in[137]),
    .X(net42));
 sky130_fd_sc_hd__clkbuf_1 input43 (.A(data_in[138]),
    .X(net43));
 sky130_fd_sc_hd__buf_1 input44 (.A(data_in[139]),
    .X(net44));
 sky130_fd_sc_hd__buf_1 input45 (.A(data_in[13]),
    .X(net45));
 sky130_fd_sc_hd__buf_1 input46 (.A(data_in[140]),
    .X(net46));
 sky130_fd_sc_hd__buf_1 input47 (.A(data_in[141]),
    .X(net47));
 sky130_fd_sc_hd__buf_1 input48 (.A(data_in[142]),
    .X(net48));
 sky130_fd_sc_hd__buf_1 input49 (.A(data_in[143]),
    .X(net49));
 sky130_fd_sc_hd__clkbuf_1 input5 (.A(data_in[103]),
    .X(net5));
 sky130_fd_sc_hd__buf_1 input50 (.A(data_in[144]),
    .X(net50));
 sky130_fd_sc_hd__buf_1 input51 (.A(data_in[145]),
    .X(net51));
 sky130_fd_sc_hd__clkbuf_2 input52 (.A(data_in[146]),
    .X(net52));
 sky130_fd_sc_hd__clkbuf_2 input53 (.A(data_in[147]),
    .X(net53));
 sky130_fd_sc_hd__clkbuf_2 input54 (.A(data_in[148]),
    .X(net54));
 sky130_fd_sc_hd__clkbuf_2 input55 (.A(data_in[149]),
    .X(net55));
 sky130_fd_sc_hd__buf_1 input56 (.A(data_in[14]),
    .X(net56));
 sky130_fd_sc_hd__clkbuf_2 input57 (.A(data_in[150]),
    .X(net57));
 sky130_fd_sc_hd__clkbuf_2 input58 (.A(data_in[151]),
    .X(net58));
 sky130_fd_sc_hd__clkbuf_2 input59 (.A(data_in[152]),
    .X(net59));
 sky130_fd_sc_hd__clkbuf_1 input6 (.A(data_in[104]),
    .X(net6));
 sky130_fd_sc_hd__buf_1 input60 (.A(data_in[153]),
    .X(net60));
 sky130_fd_sc_hd__dlymetal6s2s_1 input61 (.A(data_in[154]),
    .X(net61));
 sky130_fd_sc_hd__clkbuf_2 input62 (.A(data_in[155]),
    .X(net62));
 sky130_fd_sc_hd__clkbuf_2 input63 (.A(data_in[156]),
    .X(net63));
 sky130_fd_sc_hd__buf_1 input64 (.A(data_in[157]),
    .X(net64));
 sky130_fd_sc_hd__clkbuf_2 input65 (.A(data_in[158]),
    .X(net65));
 sky130_fd_sc_hd__clkbuf_2 input66 (.A(data_in[159]),
    .X(net66));
 sky130_fd_sc_hd__clkbuf_1 input67 (.A(data_in[15]),
    .X(net67));
 sky130_fd_sc_hd__clkbuf_2 input68 (.A(data_in[160]),
    .X(net68));
 sky130_fd_sc_hd__clkbuf_2 input69 (.A(data_in[161]),
    .X(net69));
 sky130_fd_sc_hd__buf_1 input7 (.A(data_in[105]),
    .X(net7));
 sky130_fd_sc_hd__buf_1 input70 (.A(data_in[162]),
    .X(net70));
 sky130_fd_sc_hd__clkbuf_1 input71 (.A(data_in[16]),
    .X(net71));
 sky130_fd_sc_hd__buf_1 input72 (.A(data_in[17]),
    .X(net72));
 sky130_fd_sc_hd__clkbuf_1 input73 (.A(data_in[18]),
    .X(net73));
 sky130_fd_sc_hd__clkbuf_1 input74 (.A(data_in[19]),
    .X(net74));
 sky130_fd_sc_hd__buf_1 input75 (.A(data_in[1]),
    .X(net75));
 sky130_fd_sc_hd__clkbuf_1 input76 (.A(data_in[20]),
    .X(net76));
 sky130_fd_sc_hd__clkbuf_1 input77 (.A(data_in[21]),
    .X(net77));
 sky130_fd_sc_hd__clkbuf_1 input78 (.A(data_in[22]),
    .X(net78));
 sky130_fd_sc_hd__buf_1 input79 (.A(data_in[23]),
    .X(net79));
 sky130_fd_sc_hd__buf_1 input8 (.A(data_in[106]),
    .X(net8));
 sky130_fd_sc_hd__buf_1 input80 (.A(data_in[24]),
    .X(net80));
 sky130_fd_sc_hd__buf_1 input81 (.A(data_in[25]),
    .X(net81));
 sky130_fd_sc_hd__clkbuf_1 input82 (.A(data_in[26]),
    .X(net82));
 sky130_fd_sc_hd__clkbuf_1 input83 (.A(data_in[27]),
    .X(net83));
 sky130_fd_sc_hd__clkbuf_1 input84 (.A(data_in[28]),
    .X(net84));
 sky130_fd_sc_hd__clkbuf_1 input85 (.A(data_in[29]),
    .X(net85));
 sky130_fd_sc_hd__buf_1 input86 (.A(data_in[2]),
    .X(net86));
 sky130_fd_sc_hd__clkbuf_1 input87 (.A(data_in[30]),
    .X(net87));
 sky130_fd_sc_hd__clkbuf_1 input88 (.A(data_in[31]),
    .X(net88));
 sky130_fd_sc_hd__clkbuf_1 input89 (.A(data_in[32]),
    .X(net89));
 sky130_fd_sc_hd__clkbuf_1 input9 (.A(data_in[107]),
    .X(net9));
 sky130_fd_sc_hd__clkbuf_1 input90 (.A(data_in[33]),
    .X(net90));
 sky130_fd_sc_hd__clkbuf_1 input91 (.A(data_in[34]),
    .X(net91));
 sky130_fd_sc_hd__buf_1 input92 (.A(data_in[35]),
    .X(net92));
 sky130_fd_sc_hd__clkbuf_1 input93 (.A(data_in[36]),
    .X(net93));
 sky130_fd_sc_hd__buf_1 input94 (.A(data_in[37]),
    .X(net94));
 sky130_fd_sc_hd__buf_1 input95 (.A(data_in[38]),
    .X(net95));
 sky130_fd_sc_hd__buf_1 input96 (.A(data_in[39]),
    .X(net96));
 sky130_fd_sc_hd__buf_1 input97 (.A(data_in[3]),
    .X(net97));
 sky130_fd_sc_hd__buf_1 input98 (.A(data_in[40]),
    .X(net98));
 sky130_fd_sc_hd__buf_1 input99 (.A(data_in[41]),
    .X(net99));
 sky130_fd_sc_hd__buf_12 output263 (.A(net263),
    .X(data_out[0]));
 sky130_fd_sc_hd__buf_12 output264 (.A(net264),
    .X(data_out[100]));
 sky130_fd_sc_hd__buf_12 output265 (.A(net265),
    .X(data_out[101]));
 sky130_fd_sc_hd__buf_12 output266 (.A(net266),
    .X(data_out[102]));
 sky130_fd_sc_hd__buf_12 output267 (.A(net267),
    .X(data_out[103]));
 sky130_fd_sc_hd__buf_12 output268 (.A(net268),
    .X(data_out[104]));
 sky130_fd_sc_hd__buf_12 output269 (.A(net269),
    .X(data_out[105]));
 sky130_fd_sc_hd__buf_12 output270 (.A(net270),
    .X(data_out[106]));
 sky130_fd_sc_hd__buf_12 output271 (.A(net271),
    .X(data_out[107]));
 sky130_fd_sc_hd__buf_12 output272 (.A(net272),
    .X(data_out[108]));
 sky130_fd_sc_hd__buf_12 output273 (.A(net273),
    .X(data_out[109]));
 sky130_fd_sc_hd__buf_12 output274 (.A(net274),
    .X(data_out[10]));
 sky130_fd_sc_hd__buf_12 output275 (.A(net275),
    .X(data_out[110]));
 sky130_fd_sc_hd__buf_12 output276 (.A(net276),
    .X(data_out[111]));
 sky130_fd_sc_hd__buf_12 output277 (.A(net277),
    .X(data_out[112]));
 sky130_fd_sc_hd__buf_12 output278 (.A(net278),
    .X(data_out[113]));
 sky130_fd_sc_hd__buf_12 output279 (.A(net279),
    .X(data_out[114]));
 sky130_fd_sc_hd__buf_12 output280 (.A(net280),
    .X(data_out[115]));
 sky130_fd_sc_hd__buf_12 output281 (.A(net281),
    .X(data_out[116]));
 sky130_fd_sc_hd__buf_12 output282 (.A(net282),
    .X(data_out[117]));
 sky130_fd_sc_hd__buf_12 output283 (.A(net283),
    .X(data_out[118]));
 sky130_fd_sc_hd__buf_12 output284 (.A(net284),
    .X(data_out[119]));
 sky130_fd_sc_hd__buf_12 output285 (.A(net285),
    .X(data_out[11]));
 sky130_fd_sc_hd__buf_12 output286 (.A(net286),
    .X(data_out[120]));
 sky130_fd_sc_hd__buf_12 output287 (.A(net287),
    .X(data_out[121]));
 sky130_fd_sc_hd__buf_12 output288 (.A(net288),
    .X(data_out[122]));
 sky130_fd_sc_hd__buf_12 output289 (.A(net289),
    .X(data_out[123]));
 sky130_fd_sc_hd__buf_12 output290 (.A(net290),
    .X(data_out[124]));
 sky130_fd_sc_hd__buf_12 output291 (.A(net291),
    .X(data_out[125]));
 sky130_fd_sc_hd__buf_12 output292 (.A(net292),
    .X(data_out[126]));
 sky130_fd_sc_hd__buf_12 output293 (.A(net293),
    .X(data_out[127]));
 sky130_fd_sc_hd__buf_12 output294 (.A(net294),
    .X(data_out[128]));
 sky130_fd_sc_hd__buf_12 output295 (.A(net295),
    .X(data_out[129]));
 sky130_fd_sc_hd__buf_12 output296 (.A(net296),
    .X(data_out[12]));
 sky130_fd_sc_hd__buf_12 output297 (.A(net297),
    .X(data_out[130]));
 sky130_fd_sc_hd__buf_12 output298 (.A(net298),
    .X(data_out[131]));
 sky130_fd_sc_hd__buf_12 output299 (.A(net299),
    .X(data_out[132]));
 sky130_fd_sc_hd__buf_12 output300 (.A(net300),
    .X(data_out[133]));
 sky130_fd_sc_hd__buf_12 output301 (.A(net301),
    .X(data_out[134]));
 sky130_fd_sc_hd__buf_12 output302 (.A(net302),
    .X(data_out[135]));
 sky130_fd_sc_hd__buf_12 output303 (.A(net303),
    .X(data_out[136]));
 sky130_fd_sc_hd__buf_12 output304 (.A(net304),
    .X(data_out[137]));
 sky130_fd_sc_hd__buf_12 output305 (.A(net305),
    .X(data_out[138]));
 sky130_fd_sc_hd__buf_12 output306 (.A(net306),
    .X(data_out[139]));
 sky130_fd_sc_hd__buf_12 output307 (.A(net307),
    .X(data_out[13]));
 sky130_fd_sc_hd__buf_12 output308 (.A(net308),
    .X(data_out[140]));
 sky130_fd_sc_hd__buf_12 output309 (.A(net309),
    .X(data_out[141]));
 sky130_fd_sc_hd__buf_12 output310 (.A(net310),
    .X(data_out[142]));
 sky130_fd_sc_hd__buf_12 output311 (.A(net311),
    .X(data_out[143]));
 sky130_fd_sc_hd__buf_12 output312 (.A(net312),
    .X(data_out[144]));
 sky130_fd_sc_hd__buf_12 output313 (.A(net313),
    .X(data_out[145]));
 sky130_fd_sc_hd__buf_12 output314 (.A(net314),
    .X(data_out[146]));
 sky130_fd_sc_hd__buf_12 output315 (.A(net315),
    .X(data_out[147]));
 sky130_fd_sc_hd__buf_12 output316 (.A(net316),
    .X(data_out[148]));
 sky130_fd_sc_hd__buf_12 output317 (.A(net317),
    .X(data_out[149]));
 sky130_fd_sc_hd__buf_12 output318 (.A(net318),
    .X(data_out[14]));
 sky130_fd_sc_hd__buf_12 output319 (.A(net319),
    .X(data_out[150]));
 sky130_fd_sc_hd__buf_12 output320 (.A(net320),
    .X(data_out[151]));
 sky130_fd_sc_hd__buf_12 output321 (.A(net321),
    .X(data_out[152]));
 sky130_fd_sc_hd__buf_12 output322 (.A(net322),
    .X(data_out[153]));
 sky130_fd_sc_hd__buf_12 output323 (.A(net323),
    .X(data_out[154]));
 sky130_fd_sc_hd__buf_12 output324 (.A(net324),
    .X(data_out[155]));
 sky130_fd_sc_hd__buf_12 output325 (.A(net325),
    .X(data_out[156]));
 sky130_fd_sc_hd__buf_12 output326 (.A(net326),
    .X(data_out[157]));
 sky130_fd_sc_hd__buf_12 output327 (.A(net327),
    .X(data_out[158]));
 sky130_fd_sc_hd__buf_12 output328 (.A(net328),
    .X(data_out[159]));
 sky130_fd_sc_hd__buf_12 output329 (.A(net329),
    .X(data_out[15]));
 sky130_fd_sc_hd__buf_12 output330 (.A(net330),
    .X(data_out[160]));
 sky130_fd_sc_hd__buf_12 output331 (.A(net331),
    .X(data_out[161]));
 sky130_fd_sc_hd__buf_12 output332 (.A(net332),
    .X(data_out[162]));
 sky130_fd_sc_hd__buf_12 output333 (.A(net333),
    .X(data_out[16]));
 sky130_fd_sc_hd__buf_12 output334 (.A(net334),
    .X(data_out[17]));
 sky130_fd_sc_hd__buf_12 output335 (.A(net335),
    .X(data_out[18]));
 sky130_fd_sc_hd__buf_12 output336 (.A(net336),
    .X(data_out[19]));
 sky130_fd_sc_hd__buf_12 output337 (.A(net337),
    .X(data_out[1]));
 sky130_fd_sc_hd__buf_12 output338 (.A(net338),
    .X(data_out[20]));
 sky130_fd_sc_hd__buf_12 output339 (.A(net339),
    .X(data_out[21]));
 sky130_fd_sc_hd__buf_12 output340 (.A(net340),
    .X(data_out[22]));
 sky130_fd_sc_hd__buf_12 output341 (.A(net341),
    .X(data_out[23]));
 sky130_fd_sc_hd__buf_12 output342 (.A(net342),
    .X(data_out[24]));
 sky130_fd_sc_hd__buf_12 output343 (.A(net343),
    .X(data_out[25]));
 sky130_fd_sc_hd__buf_12 output344 (.A(net344),
    .X(data_out[26]));
 sky130_fd_sc_hd__buf_12 output345 (.A(net345),
    .X(data_out[27]));
 sky130_fd_sc_hd__buf_12 output346 (.A(net346),
    .X(data_out[28]));
 sky130_fd_sc_hd__buf_12 output347 (.A(net347),
    .X(data_out[29]));
 sky130_fd_sc_hd__buf_12 output348 (.A(net348),
    .X(data_out[2]));
 sky130_fd_sc_hd__buf_12 output349 (.A(net349),
    .X(data_out[30]));
 sky130_fd_sc_hd__buf_12 output350 (.A(net350),
    .X(data_out[31]));
 sky130_fd_sc_hd__buf_12 output351 (.A(net351),
    .X(data_out[32]));
 sky130_fd_sc_hd__buf_12 output352 (.A(net352),
    .X(data_out[33]));
 sky130_fd_sc_hd__buf_12 output353 (.A(net353),
    .X(data_out[34]));
 sky130_fd_sc_hd__buf_12 output354 (.A(net354),
    .X(data_out[35]));
 sky130_fd_sc_hd__buf_12 output355 (.A(net355),
    .X(data_out[36]));
 sky130_fd_sc_hd__buf_12 output356 (.A(net356),
    .X(data_out[37]));
 sky130_fd_sc_hd__buf_12 output357 (.A(net357),
    .X(data_out[38]));
 sky130_fd_sc_hd__buf_12 output358 (.A(net358),
    .X(data_out[39]));
 sky130_fd_sc_hd__buf_12 output359 (.A(net359),
    .X(data_out[3]));
 sky130_fd_sc_hd__buf_12 output360 (.A(net360),
    .X(data_out[40]));
 sky130_fd_sc_hd__buf_12 output361 (.A(net361),
    .X(data_out[41]));
 sky130_fd_sc_hd__buf_12 output362 (.A(net362),
    .X(data_out[42]));
 sky130_fd_sc_hd__buf_12 output363 (.A(net363),
    .X(data_out[43]));
 sky130_fd_sc_hd__buf_12 output364 (.A(net364),
    .X(data_out[44]));
 sky130_fd_sc_hd__buf_12 output365 (.A(net365),
    .X(data_out[45]));
 sky130_fd_sc_hd__buf_12 output366 (.A(net366),
    .X(data_out[46]));
 sky130_fd_sc_hd__buf_12 output367 (.A(net367),
    .X(data_out[47]));
 sky130_fd_sc_hd__buf_12 output368 (.A(net368),
    .X(data_out[48]));
 sky130_fd_sc_hd__buf_12 output369 (.A(net369),
    .X(data_out[49]));
 sky130_fd_sc_hd__buf_12 output370 (.A(net370),
    .X(data_out[4]));
 sky130_fd_sc_hd__buf_12 output371 (.A(net371),
    .X(data_out[50]));
 sky130_fd_sc_hd__buf_12 output372 (.A(net372),
    .X(data_out[51]));
 sky130_fd_sc_hd__buf_12 output373 (.A(net373),
    .X(data_out[52]));
 sky130_fd_sc_hd__buf_12 output374 (.A(net374),
    .X(data_out[53]));
 sky130_fd_sc_hd__buf_12 output375 (.A(net375),
    .X(data_out[54]));
 sky130_fd_sc_hd__buf_12 output376 (.A(net376),
    .X(data_out[55]));
 sky130_fd_sc_hd__buf_12 output377 (.A(net377),
    .X(data_out[56]));
 sky130_fd_sc_hd__buf_12 output378 (.A(net378),
    .X(data_out[57]));
 sky130_fd_sc_hd__buf_12 output379 (.A(net379),
    .X(data_out[58]));
 sky130_fd_sc_hd__buf_12 output380 (.A(net380),
    .X(data_out[59]));
 sky130_fd_sc_hd__buf_12 output381 (.A(net381),
    .X(data_out[5]));
 sky130_fd_sc_hd__buf_12 output382 (.A(net382),
    .X(data_out[60]));
 sky130_fd_sc_hd__buf_12 output383 (.A(net383),
    .X(data_out[61]));
 sky130_fd_sc_hd__buf_12 output384 (.A(net384),
    .X(data_out[62]));
 sky130_fd_sc_hd__buf_12 output385 (.A(net385),
    .X(data_out[63]));
 sky130_fd_sc_hd__buf_12 output386 (.A(net386),
    .X(data_out[64]));
 sky130_fd_sc_hd__buf_12 output387 (.A(net387),
    .X(data_out[65]));
 sky130_fd_sc_hd__buf_12 output388 (.A(net388),
    .X(data_out[66]));
 sky130_fd_sc_hd__buf_12 output389 (.A(net389),
    .X(data_out[67]));
 sky130_fd_sc_hd__buf_12 output390 (.A(net390),
    .X(data_out[68]));
 sky130_fd_sc_hd__buf_12 output391 (.A(net391),
    .X(data_out[69]));
 sky130_fd_sc_hd__buf_12 output392 (.A(net392),
    .X(data_out[6]));
 sky130_fd_sc_hd__buf_12 output393 (.A(net393),
    .X(data_out[70]));
 sky130_fd_sc_hd__buf_12 output394 (.A(net394),
    .X(data_out[71]));
 sky130_fd_sc_hd__buf_12 output395 (.A(net395),
    .X(data_out[72]));
 sky130_fd_sc_hd__buf_12 output396 (.A(net396),
    .X(data_out[73]));
 sky130_fd_sc_hd__buf_12 output397 (.A(net397),
    .X(data_out[74]));
 sky130_fd_sc_hd__buf_12 output398 (.A(net398),
    .X(data_out[75]));
 sky130_fd_sc_hd__buf_12 output399 (.A(net399),
    .X(data_out[76]));
 sky130_fd_sc_hd__buf_12 output400 (.A(net400),
    .X(data_out[77]));
 sky130_fd_sc_hd__buf_12 output401 (.A(net401),
    .X(data_out[78]));
 sky130_fd_sc_hd__buf_12 output402 (.A(net402),
    .X(data_out[79]));
 sky130_fd_sc_hd__buf_12 output403 (.A(net403),
    .X(data_out[7]));
 sky130_fd_sc_hd__buf_12 output404 (.A(net404),
    .X(data_out[80]));
 sky130_fd_sc_hd__buf_12 output405 (.A(net405),
    .X(data_out[81]));
 sky130_fd_sc_hd__buf_12 output406 (.A(net406),
    .X(data_out[82]));
 sky130_fd_sc_hd__buf_12 output407 (.A(net407),
    .X(data_out[83]));
 sky130_fd_sc_hd__buf_12 output408 (.A(net408),
    .X(data_out[84]));
 sky130_fd_sc_hd__buf_12 output409 (.A(net409),
    .X(data_out[85]));
 sky130_fd_sc_hd__buf_12 output410 (.A(net410),
    .X(data_out[86]));
 sky130_fd_sc_hd__buf_12 output411 (.A(net411),
    .X(data_out[87]));
 sky130_fd_sc_hd__buf_12 output412 (.A(net412),
    .X(data_out[88]));
 sky130_fd_sc_hd__buf_12 output413 (.A(net413),
    .X(data_out[89]));
 sky130_fd_sc_hd__buf_12 output414 (.A(net414),
    .X(data_out[8]));
 sky130_fd_sc_hd__buf_12 output415 (.A(net415),
    .X(data_out[90]));
 sky130_fd_sc_hd__buf_12 output416 (.A(net416),
    .X(data_out[91]));
 sky130_fd_sc_hd__buf_12 output417 (.A(net417),
    .X(data_out[92]));
 sky130_fd_sc_hd__buf_12 output418 (.A(net418),
    .X(data_out[93]));
 sky130_fd_sc_hd__buf_12 output419 (.A(net419),
    .X(data_out[94]));
 sky130_fd_sc_hd__buf_12 output420 (.A(net420),
    .X(data_out[95]));
 sky130_fd_sc_hd__buf_12 output421 (.A(net421),
    .X(data_out[96]));
 sky130_fd_sc_hd__buf_12 output422 (.A(net422),
    .X(data_out[97]));
 sky130_fd_sc_hd__buf_12 output423 (.A(net423),
    .X(data_out[98]));
 sky130_fd_sc_hd__buf_12 output424 (.A(net424),
    .X(data_out[99]));
 sky130_fd_sc_hd__buf_12 output425 (.A(net425),
    .X(data_out[9]));
 sky130_fd_sc_hd__buf_12 output426 (.A(net426),
    .X(ki));
 sky130_fd_sc_hd__buf_12 output427 (.A(net1248),
    .X(la_data_out[100]));
 sky130_fd_sc_hd__buf_12 output428 (.A(net1249),
    .X(la_data_out[101]));
 sky130_fd_sc_hd__buf_12 output429 (.A(net1251),
    .X(la_data_out[102]));
 sky130_fd_sc_hd__buf_12 output430 (.A(net1252),
    .X(la_data_out[103]));
 sky130_fd_sc_hd__buf_12 output431 (.A(net1307),
    .X(la_data_out[104]));
 sky130_fd_sc_hd__buf_12 output432 (.A(net1253),
    .X(la_data_out[105]));
 sky130_fd_sc_hd__buf_12 output433 (.A(net1259),
    .X(la_data_out[106]));
 sky130_fd_sc_hd__buf_12 output434 (.A(net1228),
    .X(la_data_out[107]));
 sky130_fd_sc_hd__buf_12 output435 (.A(net1294),
    .X(la_data_out[108]));
 sky130_fd_sc_hd__buf_12 output436 (.A(net1256),
    .X(la_data_out[109]));
 sky130_fd_sc_hd__buf_12 output437 (.A(net1244),
    .X(la_data_out[110]));
 sky130_fd_sc_hd__buf_12 output438 (.A(net1245),
    .X(la_data_out[111]));
 sky130_fd_sc_hd__buf_12 output439 (.A(net1240),
    .X(la_data_out[112]));
 sky130_fd_sc_hd__buf_6 output440 (.A(net1359),
    .X(net1360));
 sky130_fd_sc_hd__buf_6 output441 (.A(net1425),
    .X(net1406));
 sky130_fd_sc_hd__buf_6 output442 (.A(net1423),
    .X(net1402));
 sky130_fd_sc_hd__buf_6 output443 (.A(net1429),
    .X(net1410));
 sky130_fd_sc_hd__buf_6 output444 (.A(net1427),
    .X(net1408));
 sky130_fd_sc_hd__buf_12 output445 (.A(net1238),
    .X(la_data_out[126]));
 sky130_fd_sc_hd__buf_12 output446 (.A(net1234),
    .X(la_data_out[127]));
 sky130_fd_sc_hd__buf_12 output447 (.A(net1262),
    .X(la_data_out[32]));
 sky130_fd_sc_hd__buf_12 output448 (.A(net1312),
    .X(la_data_out[33]));
 sky130_fd_sc_hd__buf_12 output449 (.A(net1260),
    .X(la_data_out[34]));
 sky130_fd_sc_hd__buf_12 output450 (.A(net1282),
    .X(la_data_out[35]));
 sky130_fd_sc_hd__buf_12 output451 (.A(net1285),
    .X(la_data_out[36]));
 sky130_fd_sc_hd__buf_12 output452 (.A(net1261),
    .X(la_data_out[37]));
 sky130_fd_sc_hd__buf_12 output453 (.A(net1315),
    .X(la_data_out[38]));
 sky130_fd_sc_hd__buf_12 output454 (.A(net1280),
    .X(la_data_out[39]));
 sky130_fd_sc_hd__buf_12 output455 (.A(net1295),
    .X(la_data_out[40]));
 sky130_fd_sc_hd__buf_12 output456 (.A(net1281),
    .X(la_data_out[41]));
 sky130_fd_sc_hd__buf_12 output457 (.A(net1284),
    .X(la_data_out[42]));
 sky130_fd_sc_hd__buf_12 output458 (.A(net1286),
    .X(la_data_out[43]));
 sky130_fd_sc_hd__buf_12 output459 (.A(net1298),
    .X(la_data_out[44]));
 sky130_fd_sc_hd__buf_12 output460 (.A(net1297),
    .X(la_data_out[45]));
 sky130_fd_sc_hd__buf_12 output461 (.A(net1265),
    .X(la_data_out[46]));
 sky130_fd_sc_hd__buf_12 output462 (.A(net1263),
    .X(la_data_out[47]));
 sky130_fd_sc_hd__buf_12 output463 (.A(net1224),
    .X(la_data_out[48]));
 sky130_fd_sc_hd__buf_12 output464 (.A(net1264),
    .X(la_data_out[49]));
 sky130_fd_sc_hd__buf_12 output465 (.A(net1227),
    .X(la_data_out[50]));
 sky130_fd_sc_hd__buf_12 output466 (.A(net1283),
    .X(la_data_out[51]));
 sky130_fd_sc_hd__buf_12 output467 (.A(net1296),
    .X(la_data_out[52]));
 sky130_fd_sc_hd__buf_12 output468 (.A(net1274),
    .X(la_data_out[53]));
 sky130_fd_sc_hd__buf_6 output469 (.A(net1399),
    .X(net1400));
 sky130_fd_sc_hd__buf_12 output470 (.A(net1273),
    .X(la_data_out[55]));
 sky130_fd_sc_hd__buf_12 output471 (.A(net1267),
    .X(la_data_out[56]));
 sky130_fd_sc_hd__buf_12 output472 (.A(net1254),
    .X(la_data_out[57]));
 sky130_fd_sc_hd__buf_12 output473 (.A(net1257),
    .X(la_data_out[58]));
 sky130_fd_sc_hd__buf_12 output474 (.A(net1271),
    .X(la_data_out[59]));
 sky130_fd_sc_hd__buf_12 output475 (.A(net1225),
    .X(la_data_out[60]));
 sky130_fd_sc_hd__buf_12 output476 (.A(net1255),
    .X(la_data_out[61]));
 sky130_fd_sc_hd__buf_12 output477 (.A(net1269),
    .X(la_data_out[62]));
 sky130_fd_sc_hd__buf_12 output478 (.A(net1272),
    .X(la_data_out[63]));
 sky130_fd_sc_hd__buf_12 output479 (.A(net1299),
    .X(la_data_out[64]));
 sky130_fd_sc_hd__buf_12 output480 (.A(net1304),
    .X(la_data_out[65]));
 sky130_fd_sc_hd__buf_12 output481 (.A(net1300),
    .X(la_data_out[66]));
 sky130_fd_sc_hd__buf_12 output482 (.A(net1305),
    .X(la_data_out[67]));
 sky130_fd_sc_hd__buf_12 output483 (.A(net1306),
    .X(la_data_out[68]));
 sky130_fd_sc_hd__buf_12 output484 (.A(net1303),
    .X(la_data_out[69]));
 sky130_fd_sc_hd__buf_12 output485 (.A(net1241),
    .X(la_data_out[70]));
 sky130_fd_sc_hd__buf_12 output486 (.A(net1242),
    .X(la_data_out[71]));
 sky130_fd_sc_hd__buf_12 output487 (.A(net1278),
    .X(la_data_out[72]));
 sky130_fd_sc_hd__buf_6 output488 (.A(net1403),
    .X(net1404));
 sky130_fd_sc_hd__buf_12 output489 (.A(net1277),
    .X(la_data_out[74]));
 sky130_fd_sc_hd__buf_12 output490 (.A(net1250),
    .X(la_data_out[75]));
 sky130_fd_sc_hd__buf_12 output491 (.A(net1275),
    .X(la_data_out[76]));
 sky130_fd_sc_hd__buf_12 output492 (.A(net1223),
    .X(la_data_out[77]));
 sky130_fd_sc_hd__buf_12 output493 (.A(net1229),
    .X(la_data_out[78]));
 sky130_fd_sc_hd__buf_12 output494 (.A(net1243),
    .X(la_data_out[79]));
 sky130_fd_sc_hd__buf_12 output495 (.A(net1236),
    .X(la_data_out[80]));
 sky130_fd_sc_hd__buf_12 output496 (.A(net1231),
    .X(la_data_out[81]));
 sky130_fd_sc_hd__buf_12 output497 (.A(net1237),
    .X(la_data_out[82]));
 sky130_fd_sc_hd__buf_12 output498 (.A(net1310),
    .X(la_data_out[83]));
 sky130_fd_sc_hd__buf_12 output499 (.A(net1309),
    .X(la_data_out[84]));
 sky130_fd_sc_hd__buf_12 output500 (.A(net1313),
    .X(la_data_out[85]));
 sky130_fd_sc_hd__buf_12 output501 (.A(net1287),
    .X(la_data_out[86]));
 sky130_fd_sc_hd__buf_12 output502 (.A(net1292),
    .X(la_data_out[87]));
 sky130_fd_sc_hd__buf_12 output503 (.A(net1289),
    .X(la_data_out[88]));
 sky130_fd_sc_hd__buf_12 output504 (.A(net1293),
    .X(la_data_out[89]));
 sky130_fd_sc_hd__buf_12 output505 (.A(net1302),
    .X(la_data_out[90]));
 sky130_fd_sc_hd__buf_12 output506 (.A(net1232),
    .X(la_data_out[91]));
 sky130_fd_sc_hd__buf_12 output507 (.A(net1233),
    .X(la_data_out[92]));
 sky130_fd_sc_hd__buf_12 output508 (.A(net1290),
    .X(la_data_out[93]));
 sky130_fd_sc_hd__buf_12 output509 (.A(net1308),
    .X(la_data_out[94]));
 sky130_fd_sc_hd__buf_12 output510 (.A(net1235),
    .X(la_data_out[95]));
 sky130_fd_sc_hd__buf_12 output511 (.A(net1301),
    .X(la_data_out[96]));
 sky130_fd_sc_hd__buf_12 output512 (.A(net1230),
    .X(la_data_out[97]));
 sky130_fd_sc_hd__buf_12 output513 (.A(net1246),
    .X(la_data_out[98]));
 sky130_fd_sc_hd__buf_12 output514 (.A(net1247),
    .X(la_data_out[99]));
 sky130_fd_sc_hd__buf_12 output515 (.A(net515),
    .X(load_data));
 sky130_fd_sc_hd__buf_12 output516 (.A(net516),
    .X(load_status[0]));
 sky130_fd_sc_hd__buf_12 output517 (.A(net517),
    .X(load_status[1]));
 sky130_fd_sc_hd__buf_12 output518 (.A(net518),
    .X(load_status[2]));
 sky130_fd_sc_hd__buf_12 output519 (.A(net519),
    .X(master_ena_proc));
 sky130_fd_sc_hd__buf_12 output520 (.A(net520),
    .X(trigLoad));
 assign la_data_out[0] = net618;
 assign la_data_out[10] = net628;
 assign la_data_out[114] = net650;
 assign la_data_out[115] = net651;
 assign la_data_out[116] = net652;
 assign la_data_out[117] = net653;
 assign la_data_out[118] = net654;
 assign la_data_out[119] = net655;
 assign la_data_out[11] = net629;
 assign la_data_out[120] = net656;
 assign la_data_out[121] = net657;
 assign la_data_out[12] = net630;
 assign la_data_out[13] = net631;
 assign la_data_out[14] = net632;
 assign la_data_out[15] = net633;
 assign la_data_out[16] = net634;
 assign la_data_out[17] = net635;
 assign la_data_out[18] = net636;
 assign la_data_out[19] = net637;
 assign la_data_out[1] = net619;
 assign la_data_out[20] = net638;
 assign la_data_out[21] = net639;
 assign la_data_out[22] = net640;
 assign la_data_out[23] = net641;
 assign la_data_out[24] = net642;
 assign la_data_out[25] = net643;
 assign la_data_out[26] = net644;
 assign la_data_out[27] = net645;
 assign la_data_out[28] = net646;
 assign la_data_out[29] = net647;
 assign la_data_out[2] = net620;
 assign la_data_out[30] = net648;
 assign la_data_out[31] = net649;
 assign la_data_out[3] = net621;
 assign la_data_out[4] = net622;
 assign la_data_out[5] = net623;
 assign la_data_out[6] = net624;
 assign la_data_out[7] = net625;
 assign la_data_out[8] = net626;
 assign la_data_out[9] = net627;
endmodule

