* NGSPICE file created from controller.ext - technology: sky130A

* Black-box entry subcircuit for sky130_fd_sc_hd__tapvpwrvgnd_1 abstract view
.subckt sky130_fd_sc_hd__tapvpwrvgnd_1 VGND VPWR
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__diode_2 abstract view
.subckt sky130_fd_sc_hd__diode_2 DIODE VGND VNB VPB VPWR
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__dfrtp_4 abstract view
.subckt sky130_fd_sc_hd__dfrtp_4 CLK D RESET_B VGND VNB VPB VPWR Q
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__inv_2 abstract view
.subckt sky130_fd_sc_hd__inv_2 A VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_ef_sc_hd__decap_12 abstract view
.subckt sky130_ef_sc_hd__decap_12 VGND VNB VPB VPWR
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__fill_1 abstract view
.subckt sky130_fd_sc_hd__fill_1 VGND VNB VPB VPWR
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__fill_2 abstract view
.subckt sky130_fd_sc_hd__fill_2 VGND VNB VPB VPWR
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__dlygate4sd3_1 abstract view
.subckt sky130_fd_sc_hd__dlygate4sd3_1 A VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__clkdlybuf4s25_1 abstract view
.subckt sky130_fd_sc_hd__clkdlybuf4s25_1 A VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__dlymetal6s2s_1 abstract view
.subckt sky130_fd_sc_hd__dlymetal6s2s_1 A VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__buf_1 abstract view
.subckt sky130_fd_sc_hd__buf_1 A VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__decap_8 abstract view
.subckt sky130_fd_sc_hd__decap_8 VGND VNB VPB VPWR
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__mux2_1 abstract view
.subckt sky130_fd_sc_hd__mux2_1 A0 A1 S VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__a311oi_1 abstract view
.subckt sky130_fd_sc_hd__a311oi_1 A1 A2 A3 B1 C1 VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__buf_12 abstract view
.subckt sky130_fd_sc_hd__buf_12 A VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__decap_6 abstract view
.subckt sky130_fd_sc_hd__decap_6 VGND VNB VPB VPWR
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__a221o_1 abstract view
.subckt sky130_fd_sc_hd__a221o_1 A1 A2 B1 B2 C1 VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__a22o_1 abstract view
.subckt sky130_fd_sc_hd__a22o_1 A1 A2 B1 B2 VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__decap_3 abstract view
.subckt sky130_fd_sc_hd__decap_3 VGND VNB VPB VPWR
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__and2_1 abstract view
.subckt sky130_fd_sc_hd__and2_1 A B VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__decap_4 abstract view
.subckt sky130_fd_sc_hd__decap_4 VGND VNB VPB VPWR
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__or4_2 abstract view
.subckt sky130_fd_sc_hd__or4_2 A B C D VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__dfrtp_1 abstract view
.subckt sky130_fd_sc_hd__dfrtp_1 CLK D RESET_B VGND VNB VPB VPWR Q
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__or4b_1 abstract view
.subckt sky130_fd_sc_hd__or4b_1 A B C D_N VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__clkbuf_16 abstract view
.subckt sky130_fd_sc_hd__clkbuf_16 A VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__dfrtp_2 abstract view
.subckt sky130_fd_sc_hd__dfrtp_2 CLK D RESET_B VGND VNB VPB VPWR Q
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__or2_2 abstract view
.subckt sky130_fd_sc_hd__or2_2 A B VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__and2_2 abstract view
.subckt sky130_fd_sc_hd__and2_2 A B VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__conb_1 abstract view
.subckt sky130_fd_sc_hd__conb_1 VGND VNB VPB VPWR HI LO
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__clkbuf_2 abstract view
.subckt sky130_fd_sc_hd__clkbuf_2 A VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__clkbuf_1 abstract view
.subckt sky130_fd_sc_hd__clkbuf_1 A VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__a311o_1 abstract view
.subckt sky130_fd_sc_hd__a311o_1 A1 A2 A3 B1 C1 VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__a211o_1 abstract view
.subckt sky130_fd_sc_hd__a211o_1 A1 A2 B1 C1 VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__nand2_1 abstract view
.subckt sky130_fd_sc_hd__nand2_1 A B VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__o2111a_1 abstract view
.subckt sky130_fd_sc_hd__o2111a_1 A1 A2 B1 C1 D1 VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__nor2_4 abstract view
.subckt sky130_fd_sc_hd__nor2_4 A B VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__nor2_1 abstract view
.subckt sky130_fd_sc_hd__nor2_1 A B VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__buf_6 abstract view
.subckt sky130_fd_sc_hd__buf_6 A VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__a21bo_1 abstract view
.subckt sky130_fd_sc_hd__a21bo_1 A1 A2 B1_N VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__a21bo_2 abstract view
.subckt sky130_fd_sc_hd__a21bo_2 A1 A2 B1_N VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__o2bb2a_1 abstract view
.subckt sky130_fd_sc_hd__o2bb2a_1 A1_N A2_N B1 B2 VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__buf_2 abstract view
.subckt sky130_fd_sc_hd__buf_2 A VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__or4bb_2 abstract view
.subckt sky130_fd_sc_hd__or4bb_2 A B C_N D_N VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__buf_8 abstract view
.subckt sky130_fd_sc_hd__buf_8 A VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__or4_1 abstract view
.subckt sky130_fd_sc_hd__or4_1 A B C D VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__or3b_1 abstract view
.subckt sky130_fd_sc_hd__or3b_1 A B C_N VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__buf_4 abstract view
.subckt sky130_fd_sc_hd__buf_4 A VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__mux2_2 abstract view
.subckt sky130_fd_sc_hd__mux2_2 A0 A1 S VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__nor4_1 abstract view
.subckt sky130_fd_sc_hd__nor4_1 A B C D VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__clkbuf_8 abstract view
.subckt sky130_fd_sc_hd__clkbuf_8 A VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__dlxtn_1 abstract view
.subckt sky130_fd_sc_hd__dlxtn_1 D GATE_N VGND VNB VPB VPWR Q
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__and3_1 abstract view
.subckt sky130_fd_sc_hd__and3_1 A B C VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__o21a_1 abstract view
.subckt sky130_fd_sc_hd__o21a_1 A1 A2 B1 VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__or3_1 abstract view
.subckt sky130_fd_sc_hd__or3_1 A B C VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__a32o_1 abstract view
.subckt sky130_fd_sc_hd__a32o_1 A1 A2 A3 B1 B2 VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__and4b_1 abstract view
.subckt sky130_fd_sc_hd__and4b_1 A_N B C D VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__a211oi_1 abstract view
.subckt sky130_fd_sc_hd__a211oi_1 A1 A2 B1 C1 VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__a211oi_4 abstract view
.subckt sky130_fd_sc_hd__a211oi_4 A1 A2 B1 C1 VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__o21ba_1 abstract view
.subckt sky130_fd_sc_hd__o21ba_1 A1 A2 B1_N VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__a32o_2 abstract view
.subckt sky130_fd_sc_hd__a32o_2 A1 A2 A3 B1 B2 VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__a21o_1 abstract view
.subckt sky130_fd_sc_hd__a21o_1 A1 A2 B1 VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__xor2_1 abstract view
.subckt sky130_fd_sc_hd__xor2_1 A B VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__or4b_2 abstract view
.subckt sky130_fd_sc_hd__or4b_2 A B C D_N VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__and4bb_2 abstract view
.subckt sky130_fd_sc_hd__and4bb_2 A_N B_N C D VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__clkbuf_4 abstract view
.subckt sky130_fd_sc_hd__clkbuf_4 A VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__nand4_1 abstract view
.subckt sky130_fd_sc_hd__nand4_1 A B C D VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__o211a_1 abstract view
.subckt sky130_fd_sc_hd__o211a_1 A1 A2 B1 C1 VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__nand2_4 abstract view
.subckt sky130_fd_sc_hd__nand2_4 A B VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__a2111o_1 abstract view
.subckt sky130_fd_sc_hd__a2111o_1 A1 A2 B1 C1 D1 VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__and4bb_1 abstract view
.subckt sky130_fd_sc_hd__and4bb_1 A_N B_N C D VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__and3b_1 abstract view
.subckt sky130_fd_sc_hd__and3b_1 A_N B C VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__and4_1 abstract view
.subckt sky130_fd_sc_hd__and4_1 A B C D VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__a41oi_1 abstract view
.subckt sky130_fd_sc_hd__a41oi_1 A1 A2 A3 A4 B1 VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__nor3_1 abstract view
.subckt sky130_fd_sc_hd__nor3_1 A B C VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__o211ai_1 abstract view
.subckt sky130_fd_sc_hd__o211ai_1 A1 A2 B1 C1 VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__and2b_1 abstract view
.subckt sky130_fd_sc_hd__and2b_1 A_N B VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__and4_2 abstract view
.subckt sky130_fd_sc_hd__and4_2 A B C D VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__a31oi_1 abstract view
.subckt sky130_fd_sc_hd__a31oi_1 A1 A2 A3 B1 VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__a31o_1 abstract view
.subckt sky130_fd_sc_hd__a31o_1 A1 A2 A3 B1 VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__a21oi_1 abstract view
.subckt sky130_fd_sc_hd__a21oi_1 A1 A2 B1 VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__and2_4 abstract view
.subckt sky130_fd_sc_hd__and2_4 A B VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__nand3_1 abstract view
.subckt sky130_fd_sc_hd__nand3_1 A B C VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__and3_4 abstract view
.subckt sky130_fd_sc_hd__and3_4 A B C VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__nand2_2 abstract view
.subckt sky130_fd_sc_hd__nand2_2 A B VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__nor2_2 abstract view
.subckt sky130_fd_sc_hd__nor2_2 A B VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__or2_1 abstract view
.subckt sky130_fd_sc_hd__or2_1 A B VGND VNB VPB VPWR X
.ends

.subckt controller becStatus[0] becStatus[1] becStatus[2] becStatus[3] data_in[0]
+ data_in[100] data_in[101] data_in[102] data_in[103] data_in[104] data_in[105] data_in[106]
+ data_in[107] data_in[108] data_in[109] data_in[10] data_in[110] data_in[111] data_in[112]
+ data_in[113] data_in[114] data_in[115] data_in[116] data_in[117] data_in[118] data_in[119]
+ data_in[11] data_in[120] data_in[121] data_in[122] data_in[123] data_in[124] data_in[125]
+ data_in[126] data_in[127] data_in[128] data_in[129] data_in[12] data_in[130] data_in[131]
+ data_in[132] data_in[133] data_in[134] data_in[135] data_in[136] data_in[137] data_in[138]
+ data_in[139] data_in[13] data_in[140] data_in[141] data_in[142] data_in[143] data_in[144]
+ data_in[145] data_in[146] data_in[147] data_in[148] data_in[149] data_in[14] data_in[150]
+ data_in[151] data_in[152] data_in[153] data_in[154] data_in[155] data_in[156] data_in[157]
+ data_in[158] data_in[159] data_in[15] data_in[160] data_in[161] data_in[162] data_in[16]
+ data_in[17] data_in[18] data_in[19] data_in[1] data_in[20] data_in[21] data_in[22]
+ data_in[23] data_in[24] data_in[25] data_in[26] data_in[27] data_in[28] data_in[29]
+ data_in[2] data_in[30] data_in[31] data_in[32] data_in[33] data_in[34] data_in[35]
+ data_in[36] data_in[37] data_in[38] data_in[39] data_in[3] data_in[40] data_in[41]
+ data_in[42] data_in[43] data_in[44] data_in[45] data_in[46] data_in[47] data_in[48]
+ data_in[49] data_in[4] data_in[50] data_in[51] data_in[52] data_in[53] data_in[54]
+ data_in[55] data_in[56] data_in[57] data_in[58] data_in[59] data_in[5] data_in[60]
+ data_in[61] data_in[62] data_in[63] data_in[64] data_in[65] data_in[66] data_in[67]
+ data_in[68] data_in[69] data_in[6] data_in[70] data_in[71] data_in[72] data_in[73]
+ data_in[74] data_in[75] data_in[76] data_in[77] data_in[78] data_in[79] data_in[7]
+ data_in[80] data_in[81] data_in[82] data_in[83] data_in[84] data_in[85] data_in[86]
+ data_in[87] data_in[88] data_in[89] data_in[8] data_in[90] data_in[91] data_in[92]
+ data_in[93] data_in[94] data_in[95] data_in[96] data_in[97] data_in[98] data_in[99]
+ data_in[9] data_out[0] data_out[100] data_out[101] data_out[102] data_out[103] data_out[104]
+ data_out[105] data_out[106] data_out[107] data_out[108] data_out[109] data_out[10]
+ data_out[110] data_out[111] data_out[112] data_out[113] data_out[114] data_out[115]
+ data_out[116] data_out[117] data_out[118] data_out[119] data_out[11] data_out[120]
+ data_out[121] data_out[122] data_out[123] data_out[124] data_out[125] data_out[126]
+ data_out[127] data_out[128] data_out[129] data_out[12] data_out[130] data_out[131]
+ data_out[132] data_out[133] data_out[134] data_out[135] data_out[136] data_out[137]
+ data_out[138] data_out[139] data_out[13] data_out[140] data_out[141] data_out[142]
+ data_out[143] data_out[144] data_out[145] data_out[146] data_out[147] data_out[148]
+ data_out[149] data_out[14] data_out[150] data_out[151] data_out[152] data_out[153]
+ data_out[154] data_out[155] data_out[156] data_out[157] data_out[158] data_out[159]
+ data_out[15] data_out[160] data_out[161] data_out[162] data_out[16] data_out[17]
+ data_out[18] data_out[19] data_out[1] data_out[20] data_out[21] data_out[22] data_out[23]
+ data_out[24] data_out[25] data_out[26] data_out[27] data_out[28] data_out[29] data_out[2]
+ data_out[30] data_out[31] data_out[32] data_out[33] data_out[34] data_out[35] data_out[36]
+ data_out[37] data_out[38] data_out[39] data_out[3] data_out[40] data_out[41] data_out[42]
+ data_out[43] data_out[44] data_out[45] data_out[46] data_out[47] data_out[48] data_out[49]
+ data_out[4] data_out[50] data_out[51] data_out[52] data_out[53] data_out[54] data_out[55]
+ data_out[56] data_out[57] data_out[58] data_out[59] data_out[5] data_out[60] data_out[61]
+ data_out[62] data_out[63] data_out[64] data_out[65] data_out[66] data_out[67] data_out[68]
+ data_out[69] data_out[6] data_out[70] data_out[71] data_out[72] data_out[73] data_out[74]
+ data_out[75] data_out[76] data_out[77] data_out[78] data_out[79] data_out[7] data_out[80]
+ data_out[81] data_out[82] data_out[83] data_out[84] data_out[85] data_out[86] data_out[87]
+ data_out[88] data_out[89] data_out[8] data_out[90] data_out[91] data_out[92] data_out[93]
+ data_out[94] data_out[95] data_out[96] data_out[97] data_out[98] data_out[99] data_out[9]
+ ki la_data_in[0] la_data_in[100] la_data_in[101] la_data_in[102] la_data_in[103]
+ la_data_in[104] la_data_in[105] la_data_in[106] la_data_in[107] la_data_in[108]
+ la_data_in[109] la_data_in[10] la_data_in[110] la_data_in[111] la_data_in[112] la_data_in[113]
+ la_data_in[114] la_data_in[115] la_data_in[116] la_data_in[117] la_data_in[118]
+ la_data_in[119] la_data_in[11] la_data_in[120] la_data_in[121] la_data_in[122] la_data_in[123]
+ la_data_in[124] la_data_in[125] la_data_in[126] la_data_in[127] la_data_in[12] la_data_in[13]
+ la_data_in[14] la_data_in[15] la_data_in[16] la_data_in[17] la_data_in[18] la_data_in[19]
+ la_data_in[1] la_data_in[20] la_data_in[21] la_data_in[22] la_data_in[23] la_data_in[24]
+ la_data_in[25] la_data_in[26] la_data_in[27] la_data_in[28] la_data_in[29] la_data_in[2]
+ la_data_in[30] la_data_in[31] la_data_in[32] la_data_in[33] la_data_in[34] la_data_in[35]
+ la_data_in[36] la_data_in[37] la_data_in[38] la_data_in[39] la_data_in[3] la_data_in[40]
+ la_data_in[41] la_data_in[42] la_data_in[43] la_data_in[44] la_data_in[45] la_data_in[46]
+ la_data_in[47] la_data_in[48] la_data_in[49] la_data_in[4] la_data_in[50] la_data_in[51]
+ la_data_in[52] la_data_in[53] la_data_in[54] la_data_in[55] la_data_in[56] la_data_in[57]
+ la_data_in[58] la_data_in[59] la_data_in[5] la_data_in[60] la_data_in[61] la_data_in[62]
+ la_data_in[63] la_data_in[64] la_data_in[65] la_data_in[66] la_data_in[67] la_data_in[68]
+ la_data_in[69] la_data_in[6] la_data_in[70] la_data_in[71] la_data_in[72] la_data_in[73]
+ la_data_in[74] la_data_in[75] la_data_in[76] la_data_in[77] la_data_in[78] la_data_in[79]
+ la_data_in[7] la_data_in[80] la_data_in[81] la_data_in[82] la_data_in[83] la_data_in[84]
+ la_data_in[85] la_data_in[86] la_data_in[87] la_data_in[88] la_data_in[89] la_data_in[8]
+ la_data_in[90] la_data_in[91] la_data_in[92] la_data_in[93] la_data_in[94] la_data_in[95]
+ la_data_in[96] la_data_in[97] la_data_in[98] la_data_in[99] la_data_in[9] la_data_out[0]
+ la_data_out[100] la_data_out[101] la_data_out[102] la_data_out[103] la_data_out[104]
+ la_data_out[105] la_data_out[106] la_data_out[107] la_data_out[108] la_data_out[109]
+ la_data_out[10] la_data_out[110] la_data_out[111] la_data_out[112] la_data_out[113]
+ la_data_out[114] la_data_out[115] la_data_out[116] la_data_out[117] la_data_out[118]
+ la_data_out[119] la_data_out[11] la_data_out[120] la_data_out[121] la_data_out[122]
+ la_data_out[123] la_data_out[124] la_data_out[125] la_data_out[126] la_data_out[127]
+ la_data_out[12] la_data_out[13] la_data_out[14] la_data_out[15] la_data_out[16]
+ la_data_out[17] la_data_out[18] la_data_out[19] la_data_out[1] la_data_out[20] la_data_out[21]
+ la_data_out[22] la_data_out[23] la_data_out[24] la_data_out[25] la_data_out[26]
+ la_data_out[27] la_data_out[28] la_data_out[29] la_data_out[2] la_data_out[30] la_data_out[31]
+ la_data_out[32] la_data_out[33] la_data_out[34] la_data_out[35] la_data_out[36]
+ la_data_out[37] la_data_out[38] la_data_out[39] la_data_out[3] la_data_out[40] la_data_out[41]
+ la_data_out[42] la_data_out[43] la_data_out[44] la_data_out[45] la_data_out[46]
+ la_data_out[47] la_data_out[48] la_data_out[49] la_data_out[4] la_data_out[50] la_data_out[51]
+ la_data_out[52] la_data_out[53] la_data_out[54] la_data_out[55] la_data_out[56]
+ la_data_out[57] la_data_out[58] la_data_out[59] la_data_out[5] la_data_out[60] la_data_out[61]
+ la_data_out[62] la_data_out[63] la_data_out[64] la_data_out[65] la_data_out[66]
+ la_data_out[67] la_data_out[68] la_data_out[69] la_data_out[6] la_data_out[70] la_data_out[71]
+ la_data_out[72] la_data_out[73] la_data_out[74] la_data_out[75] la_data_out[76]
+ la_data_out[77] la_data_out[78] la_data_out[79] la_data_out[7] la_data_out[80] la_data_out[81]
+ la_data_out[82] la_data_out[83] la_data_out[84] la_data_out[85] la_data_out[86]
+ la_data_out[87] la_data_out[88] la_data_out[89] la_data_out[8] la_data_out[90] la_data_out[91]
+ la_data_out[92] la_data_out[93] la_data_out[94] la_data_out[95] la_data_out[96]
+ la_data_out[97] la_data_out[98] la_data_out[99] la_data_out[9] la_oenb[0] la_oenb[100]
+ la_oenb[101] la_oenb[102] la_oenb[103] la_oenb[104] la_oenb[105] la_oenb[106] la_oenb[107]
+ la_oenb[108] la_oenb[109] la_oenb[10] la_oenb[110] la_oenb[111] la_oenb[112] la_oenb[113]
+ la_oenb[114] la_oenb[115] la_oenb[116] la_oenb[117] la_oenb[118] la_oenb[119] la_oenb[11]
+ la_oenb[120] la_oenb[121] la_oenb[122] la_oenb[123] la_oenb[124] la_oenb[125] la_oenb[126]
+ la_oenb[127] la_oenb[12] la_oenb[13] la_oenb[14] la_oenb[15] la_oenb[16] la_oenb[17]
+ la_oenb[18] la_oenb[19] la_oenb[1] la_oenb[20] la_oenb[21] la_oenb[22] la_oenb[23]
+ la_oenb[24] la_oenb[25] la_oenb[26] la_oenb[27] la_oenb[28] la_oenb[29] la_oenb[2]
+ la_oenb[30] la_oenb[31] la_oenb[32] la_oenb[33] la_oenb[34] la_oenb[35] la_oenb[36]
+ la_oenb[37] la_oenb[38] la_oenb[39] la_oenb[3] la_oenb[40] la_oenb[41] la_oenb[42]
+ la_oenb[43] la_oenb[44] la_oenb[45] la_oenb[46] la_oenb[47] la_oenb[48] la_oenb[49]
+ la_oenb[4] la_oenb[50] la_oenb[51] la_oenb[52] la_oenb[53] la_oenb[54] la_oenb[55]
+ la_oenb[56] la_oenb[57] la_oenb[58] la_oenb[59] la_oenb[5] la_oenb[60] la_oenb[61]
+ la_oenb[62] la_oenb[63] la_oenb[64] la_oenb[65] la_oenb[66] la_oenb[67] la_oenb[68]
+ la_oenb[69] la_oenb[6] la_oenb[70] la_oenb[71] la_oenb[72] la_oenb[73] la_oenb[74]
+ la_oenb[75] la_oenb[76] la_oenb[77] la_oenb[78] la_oenb[79] la_oenb[7] la_oenb[80]
+ la_oenb[81] la_oenb[82] la_oenb[83] la_oenb[84] la_oenb[85] la_oenb[86] la_oenb[87]
+ la_oenb[88] la_oenb[89] la_oenb[8] la_oenb[90] la_oenb[91] la_oenb[92] la_oenb[93]
+ la_oenb[94] la_oenb[95] la_oenb[96] la_oenb[97] la_oenb[98] la_oenb[99] la_oenb[9]
+ load_data load_status[0] load_status[1] load_status[2] master_ena_proc next_key
+ slv_done trigLoad vccd1 vssd1 wb_clk_i wb_rst_i
XTAP_199 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_188 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_177 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__1151__B1 _1183_/B1 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_2106_ _2106_/CLK _2106_/D _1849_/Y vssd1 vssd1 vccd1 vccd1 _2106_/Q sky130_fd_sc_hd__dfrtp_4
X_2037_ _2065_/A vssd1 vssd1 vccd1 vccd1 _2037_/Y sky130_fd_sc_hd__inv_2
XFILLER_0_18_701 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_45_531 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_17_200 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_17_222 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_45_553 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_17_255 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__1206__A1 input70/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_32_203 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__1509__A2 _1519_/A2 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xhold351 hold365/X vssd1 vssd1 vccd1 vccd1 hold351/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold362 la_data_in[72] vssd1 vssd1 vccd1 vccd1 hold362/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold340 _1274_/X vssd1 vssd1 vccd1 vccd1 hold340/X sky130_fd_sc_hd__clkdlybuf4s25_1
Xhold395 la_data_in[67] vssd1 vssd1 vccd1 vccd1 hold395/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold373 _1262_/X vssd1 vssd1 vccd1 vccd1 hold373/X sky130_fd_sc_hd__dlymetal6s2s_1
Xhold384 _1232_/X vssd1 vssd1 vccd1 vccd1 hold384/X sky130_fd_sc_hd__buf_1
XANTENNA__1142__A0 _2185_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_3_609 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_36_597 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_23_236 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_23_269 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_48_15 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_48_48 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_48_37 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_48_26 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_1270_ _1269_/X _2221_/Q _1318_/S vssd1 vssd1 vccd1 vccd1 _1270_/X sky130_fd_sc_hd__mux2_1
XANTENNA__1133__B1 _1157_/B1 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_6_425 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_54_361 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_42_523 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_0985_ _0971_/C hold428/X _0983_/B hold36/X _0973_/B vssd1 vssd1 vccd1 vccd1 _0985_/Y
+ sky130_fd_sc_hd__a311oi_1
XFILLER_0_14_214 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
Xoutput401 _1720_/X vssd1 vssd1 vccd1 vccd1 data_out[78] sky130_fd_sc_hd__buf_12
XFILLER_0_42_578 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_30_707 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
Xoutput412 _1730_/X vssd1 vssd1 vccd1 vccd1 data_out[88] sky130_fd_sc_hd__buf_12
Xoutput423 _1740_/X vssd1 vssd1 vccd1 vccd1 data_out[98] sky130_fd_sc_hd__buf_12
Xoutput434 hold571/X vssd1 vssd1 vccd1 vccd1 la_data_out[107] sky130_fd_sc_hd__buf_12
X_1606_ hold220/X hold972/X _1632_/S vssd1 vssd1 vccd1 vccd1 _2083_/D sky130_fd_sc_hd__mux2_1
Xoutput445 hold581/X vssd1 vssd1 vccd1 vccd1 la_data_out[126] sky130_fd_sc_hd__buf_12
Xoutput478 hold615/X vssd1 vssd1 vccd1 vccd1 la_data_out[63] sky130_fd_sc_hd__buf_12
Xoutput467 hold639/X vssd1 vssd1 vccd1 vccd1 la_data_out[52] sky130_fd_sc_hd__buf_12
Xoutput456 hold624/X vssd1 vssd1 vccd1 vccd1 la_data_out[41] sky130_fd_sc_hd__buf_12
XFILLER_0_10_475 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xoutput489 hold620/X vssd1 vssd1 vccd1 vccd1 la_data_out[74] sky130_fd_sc_hd__buf_12
X_1537_ _1537_/A1 _1197_/D _1541_/B1 _2118_/Q hold95/X vssd1 vssd1 vccd1 vccd1 _1537_/X
+ sky130_fd_sc_hd__a221o_1
X_1468_ _1310_/A hold6/X _1541_/B1 _2162_/Q vssd1 vssd1 vccd1 vccd1 hold7/A sky130_fd_sc_hd__a22o_1
XANTENNA__1124__A0 _2194_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_1399_ _1398_/X hold775/X _1435_/S vssd1 vssd1 vccd1 vccd1 _2178_/D sky130_fd_sc_hd__mux2_1
XFILLER_0_54_80 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_49_111 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA_fanout544_A _1641_/Y vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_49_166 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_52_309 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_18_531 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_45_361 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_18_575 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xhold170 _1473_/X vssd1 vssd1 vccd1 vccd1 hold170/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold181 hold210/X vssd1 vssd1 vccd1 vccd1 hold181/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold192 _1551_/X vssd1 vssd1 vccd1 vccd1 hold192/X sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_18_29 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__1115__B1 _1183_/B1 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_hold923_A _2177_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_55_158 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_50_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_55_169 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_24_523 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_24_545 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_24_589 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_11_228 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_1322_ _1349_/A _1322_/B vssd1 vssd1 vccd1 vccd1 _1322_/X sky130_fd_sc_hd__and2_1
X_1253_ _1271_/A _1253_/B vssd1 vssd1 vccd1 vccd1 _1253_/X sky130_fd_sc_hd__and2_1
XANTENNA__1902__A _1913_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_1184_ _2164_/Q _2072_/Q _1188_/S vssd1 vssd1 vccd1 vccd1 _1184_/X sky130_fd_sc_hd__mux2_1
XANTENNA_clkbuf_leaf_4_wb_clk_i_A clkbuf_leaf_9_wb_clk_i/A vssd1 vssd1 vccd1 vccd1
+ sky130_fd_sc_hd__diode_2
XFILLER_0_46_103 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_19_317 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_24_83 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_46_136 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_0968_ _0977_/C _0978_/A _0978_/B _0973_/D vssd1 vssd1 vccd1 vccd1 _0969_/C sky130_fd_sc_hd__or4_2
XFILLER_0_6_288 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_40_93 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__1593__B1 _1623_/B1 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_30_515 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
Xoutput275 _1752_/X vssd1 vssd1 vccd1 vccd1 data_out[110] sky130_fd_sc_hd__buf_12
Xoutput264 _1742_/X vssd1 vssd1 vccd1 vccd1 data_out[100] sky130_fd_sc_hd__buf_12
Xoutput286 _1762_/X vssd1 vssd1 vccd1 vccd1 data_out[120] sky130_fd_sc_hd__buf_12
XFILLER_0_10_250 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
Xoutput297 _1772_/X vssd1 vssd1 vccd1 vccd1 data_out[130] sky130_fd_sc_hd__buf_12
XANTENNA__1812__A _2070_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_18_361 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_37_169 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_18_372 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_33_386 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__1706__B _1715_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_1940_ _1941_/A vssd1 vssd1 vccd1 vccd1 _1940_/Y sky130_fd_sc_hd__inv_2
X_1871_ _2002_/A vssd1 vssd1 vccd1 vccd1 _1871_/Y sky130_fd_sc_hd__inv_2
XFILLER_0_28_158 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_37_670 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_51_161 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
Xhold906 _2153_/Q vssd1 vssd1 vccd1 vccd1 hold906/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold917 la_data_in[7] vssd1 vssd1 vccd1 vccd1 hold917/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold928 _1584_/X vssd1 vssd1 vccd1 vccd1 _2094_/D sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_51_194 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
Xhold939 _1580_/X vssd1 vssd1 vccd1 vccd1 _2096_/D sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA__1108__S _1188_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_1305_ input33/X _1527_/A2 _1541_/B1 _2210_/Q hold95/X vssd1 vssd1 vccd1 vccd1 hold96/A
+ sky130_fd_sc_hd__a221o_1
X_2285_ _2312_/CLK _2285_/D _2024_/Y vssd1 vssd1 vccd1 vccd1 _2285_/Q sky130_fd_sc_hd__dfrtp_1
X_1236_ input59/X _1495_/A2 _1495_/B1 _2233_/Q hold410/X vssd1 vssd1 vccd1 vccd1 _1236_/X
+ sky130_fd_sc_hd__a221o_1
X_1167_ hold629/X _1183_/A2 _1183_/B1 _1166_/X vssd1 vssd1 vccd1 vccd1 _2261_/D sky130_fd_sc_hd__a22o_1
XFILLER_0_19_103 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_1098_ _2207_/Q _2115_/Q _1112_/S vssd1 vssd1 vccd1 vccd1 _1098_/X sky130_fd_sc_hd__mux2_1
XFILLER_0_47_456 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_47_467 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_19_169 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_34_117 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_43_640 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__1097__A2 _1097_/A2 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_38_489 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_25_128 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XANTENNA_hold990_A _2093_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_34_662 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_33_150 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_34_673 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XANTENNA__1557__B1 _1623_/B1 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_21_323 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_21_345 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_33_183 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_21_389 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_507 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_518 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_529 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_56_15 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_2070_ _2164_/CLK hold51/X _0956_/Y vssd1 vssd1 vccd1 vccd1 _2070_/Q sky130_fd_sc_hd__dfrtp_4
X_1021_ hold38/X _1194_/A _1191_/B hold430/X vssd1 vssd1 vccd1 vccd1 _1021_/X sky130_fd_sc_hd__or4b_1
XFILLER_0_8_317 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_56_253 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_1923_ _1941_/A vssd1 vssd1 vccd1 vccd1 _1923_/Y sky130_fd_sc_hd__inv_2
XFILLER_0_29_489 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XANTENNA__1260__A2 _1519_/A2 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_1854_ _1988_/A vssd1 vssd1 vccd1 vccd1 _1854_/Y sky130_fd_sc_hd__inv_2
X_1785_ _2223_/Q _1798_/B vssd1 vssd1 vccd1 vccd1 _1785_/X sky130_fd_sc_hd__and2_1
XFILLER_0_12_301 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
Xhold703 hold703/A vssd1 vssd1 vccd1 vccd1 la_data_out[113] sky130_fd_sc_hd__buf_12
XFILLER_0_25_673 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
Xhold736 hold861/X vssd1 vssd1 vccd1 vccd1 hold736/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold714 hold906/X vssd1 vssd1 vccd1 vccd1 hold714/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold725 hold877/X vssd1 vssd1 vccd1 vccd1 hold725/X sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_12_356 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
Xhold769 _2160_/Q vssd1 vssd1 vccd1 vccd1 hold769/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold747 hold747/A vssd1 vssd1 vccd1 vccd1 la_data_out[73] sky130_fd_sc_hd__buf_12
Xhold758 hold785/X vssd1 vssd1 vccd1 vccd1 hold758/X sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_34_3 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_2268_ _2300_/CLK _2268_/D _2007_/Y vssd1 vssd1 vccd1 vccd1 _2268_/Q sky130_fd_sc_hd__dfrtp_1
X_1219_ hold416/X _2238_/Q _1252_/S vssd1 vssd1 vccd1 vccd1 _1219_/X sky130_fd_sc_hd__mux2_1
XANTENNA__1079__A2 _1095_/A2 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_2199_ _2219_/CLK _2199_/D _1939_/Y vssd1 vssd1 vccd1 vccd1 _2199_/Q sky130_fd_sc_hd__dfrtp_4
XFILLER_0_48_710 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_7_383 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_16_651 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_50_429 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_16_684 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__1539__B1 _1541_/B1 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_43_492 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_31_665 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_30_197 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xhold30 hold30/A vssd1 vssd1 vccd1 vccd1 hold30/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold41 hold41/A vssd1 vssd1 vccd1 vccd1 hold41/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold63 hold63/A vssd1 vssd1 vccd1 vccd1 hold63/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold52 hold52/A vssd1 vssd1 vccd1 vccd1 hold52/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold74 hold74/A vssd1 vssd1 vccd1 vccd1 hold74/X sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_26_29 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
Xhold85 hold85/A vssd1 vssd1 vccd1 vccd1 hold85/X sky130_fd_sc_hd__buf_1
Xhold96 hold96/A vssd1 vssd1 vccd1 vccd1 hold96/X sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_38_220 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_54_713 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__1227__C1 hold422/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_53_212 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_26_448 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_53_245 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_53_234 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
Xclkbuf_leaf_14_wb_clk_i clkbuf_1_1__f_wb_clk_i/X vssd1 vssd1 vccd1 vccd1 _2239_/CLK
+ sky130_fd_sc_hd__clkbuf_16
XFILLER_0_41_429 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_1570_ hold245/X hold937/X hold81/X vssd1 vssd1 vccd1 vccd1 _2101_/D sky130_fd_sc_hd__mux2_1
XANTENNA_5 la_data_in[32] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_22_665 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_315 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_304 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_326 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_337 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_348 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_359 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_2122_ _2219_/CLK _2122_/D _1865_/Y vssd1 vssd1 vccd1 vccd1 _2122_/Q sky130_fd_sc_hd__dfrtp_2
X_2053_ _2065_/A vssd1 vssd1 vccd1 vccd1 _2053_/Y sky130_fd_sc_hd__inv_2
X_1004_ _2248_/Q _1445_/A vssd1 vssd1 vccd1 vccd1 _1805_/A sky130_fd_sc_hd__or2_2
XANTENNA__1481__A2 _1503_/A2 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_45_713 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_29_253 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__1218__C1 hold415/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_17_415 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_29_297 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__1233__A2 _1503_/A2 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_1906_ _1916_/A vssd1 vssd1 vccd1 vccd1 _1906_/Y sky130_fd_sc_hd__inv_2
X_1837_ _1852_/A vssd1 vssd1 vccd1 vccd1 _1837_/Y sky130_fd_sc_hd__inv_2
Xhold511 _1810_/B vssd1 vssd1 vccd1 vccd1 _1397_/B sky130_fd_sc_hd__dlygate4sd3_1
Xhold500 _1265_/X vssd1 vssd1 vccd1 vccd1 hold500/X sky130_fd_sc_hd__buf_1
Xhold522 _1386_/X vssd1 vssd1 vccd1 vccd1 hold522/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold533 la_data_in[22] vssd1 vssd1 vccd1 vccd1 hold533/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold544 _1449_/X vssd1 vssd1 vccd1 vccd1 _2160_/D sky130_fd_sc_hd__dlygate4sd3_1
X_1768_ _2206_/Q _1804_/B vssd1 vssd1 vccd1 vccd1 _1768_/X sky130_fd_sc_hd__and2_2
X_1699_ _2127_/Q _1715_/B vssd1 vssd1 vccd1 vccd1 _1699_/X sky130_fd_sc_hd__and2_1
XFILLER_0_12_197 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xhold555 _1192_/X vssd1 vssd1 vccd1 vccd1 _1194_/B sky130_fd_sc_hd__dlygate4sd3_1
Xhold588 hold670/X vssd1 vssd1 vccd1 vccd1 hold588/X sky130_fd_sc_hd__dlymetal6s2s_1
Xhold577 hold714/X vssd1 vssd1 vccd1 vccd1 hold577/X sky130_fd_sc_hd__dlymetal6s2s_1
Xhold566 hold677/X vssd1 vssd1 vccd1 vccd1 hold566/X sky130_fd_sc_hd__dlymetal6s2s_1
Xhold599 hold732/X vssd1 vssd1 vccd1 vccd1 hold599/X sky130_fd_sc_hd__dlymetal6s2s_1
XFILLER_0_0_592 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_871 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_860 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_fanout574_A _1569_/B1 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_893 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_882 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_57_91 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__1457__C1 _1545_/B1 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_36_713 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__1224__A2 _1503_/A2 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xcontroller_630 vssd1 vssd1 vccd1 vccd1 controller_630/HI la_data_out[12] sky130_fd_sc_hd__conb_1
Xcontroller_641 vssd1 vssd1 vccd1 vccd1 controller_641/HI la_data_out[23] sky130_fd_sc_hd__conb_1
Xcontroller_652 vssd1 vssd1 vccd1 vccd1 controller_652/HI la_data_out[116] sky130_fd_sc_hd__conb_1
XANTENNA_hold786_A _2109_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_31_462 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_31_484 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA_hold953_A _2175_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xinput120 data_in[60] vssd1 vssd1 vccd1 vccd1 _1511_/A1 sky130_fd_sc_hd__dlymetal6s2s_1
Xinput142 data_in[80] vssd1 vssd1 vccd1 vccd1 _1471_/A1 sky130_fd_sc_hd__dlymetal6s2s_1
Xinput131 data_in[70] vssd1 vssd1 vccd1 vccd1 _1491_/A1 sky130_fd_sc_hd__clkbuf_2
Xinput153 data_in[90] vssd1 vssd1 vccd1 vccd1 _1422_/A1 sky130_fd_sc_hd__buf_1
Xinput164 hold47/X vssd1 vssd1 vccd1 vccd1 hold48/A sky130_fd_sc_hd__clkbuf_1
Xinput186 hold15/X vssd1 vssd1 vccd1 vccd1 hold16/A sky130_fd_sc_hd__clkbuf_1
Xinput175 hold29/X vssd1 vssd1 vccd1 vccd1 hold30/A sky130_fd_sc_hd__clkbuf_1
XANTENNA__1160__A1 _2084_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__1730__A _2168_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xinput197 hold174/X vssd1 vssd1 vccd1 vccd1 hold175/A sky130_fd_sc_hd__clkbuf_1
XFILLER_0_39_551 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_1622_ _1621_/X hold958/X _1622_/S vssd1 vssd1 vccd1 vccd1 _2075_/D sky130_fd_sc_hd__mux2_1
XFILLER_0_22_462 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__1905__A _1913_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_1553_ input96/X _1637_/B _1635_/C _2110_/Q hold254/X vssd1 vssd1 vccd1 vccd1 _1553_/X
+ sky130_fd_sc_hd__a221o_1
X_1484_ _1483_/X _2144_/Q _1504_/S vssd1 vssd1 vccd1 vccd1 _1484_/X sky130_fd_sc_hd__mux2_1
XTAP_123 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_1_378 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_1_389 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_145 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_134 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_156 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_189 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_178 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_167 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_27_72 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_2105_ _2168_/CLK _2105_/D _1848_/Y vssd1 vssd1 vccd1 vccd1 _2105_/Q sky130_fd_sc_hd__dfrtp_4
X_2036_ _2065_/A vssd1 vssd1 vccd1 vccd1 _2036_/Y sky130_fd_sc_hd__inv_2
XFILLER_0_49_337 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_9_401 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_45_521 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_17_212 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_18_713 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__1206__A2 _1197_/D vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_45_598 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_45_587 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xhold341 _1275_/X vssd1 vssd1 vccd1 vccd1 hold341/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold352 hold352/A vssd1 vssd1 vccd1 vccd1 _1286_/B sky130_fd_sc_hd__dlygate4sd3_1
Xhold330 la_data_in[66] vssd1 vssd1 vccd1 vccd1 hold330/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold374 _1263_/X vssd1 vssd1 vccd1 vccd1 hold374/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold385 _1489_/X vssd1 vssd1 vccd1 vccd1 hold385/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold363 _1231_/X vssd1 vssd1 vccd1 vccd1 _2234_/D sky130_fd_sc_hd__dlygate4sd3_1
Xhold396 _1246_/X vssd1 vssd1 vccd1 vccd1 _2229_/D sky130_fd_sc_hd__dlygate4sd3_1
XTAP_690 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__1142__A1 _2093_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_36_510 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_51_502 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_36_587 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__1725__A _2163_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_27_521 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_39_381 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_13_63 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_54_373 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_0984_ _0971_/C hold428/X _0983_/B hold36/X _0973_/B vssd1 vssd1 vccd1 vccd1 hold37/A
+ sky130_fd_sc_hd__a311o_1
XFILLER_0_14_226 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xoutput402 _1721_/X vssd1 vssd1 vccd1 vccd1 data_out[79] sky130_fd_sc_hd__buf_12
XFILLER_0_42_568 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xoutput413 _1731_/X vssd1 vssd1 vccd1 vccd1 data_out[89] sky130_fd_sc_hd__buf_12
Xoutput424 _1741_/X vssd1 vssd1 vccd1 vccd1 data_out[99] sky130_fd_sc_hd__buf_12
Xoutput435 hold637/X vssd1 vssd1 vccd1 vccd1 la_data_out[108] sky130_fd_sc_hd__buf_12
X_1605_ input45/X _1623_/A2 _1623_/B1 _2084_/Q hold219/X vssd1 vssd1 vccd1 vccd1 _1605_/X
+ sky130_fd_sc_hd__a221o_1
Xoutput446 hold577/X vssd1 vssd1 vccd1 vccd1 la_data_out[127] sky130_fd_sc_hd__buf_12
Xoutput468 hold617/X vssd1 vssd1 vccd1 vccd1 la_data_out[53] sky130_fd_sc_hd__buf_12
Xoutput457 hold627/X vssd1 vssd1 vccd1 vccd1 la_data_out[42] sky130_fd_sc_hd__buf_12
X_1536_ _1535_/X _2118_/Q hold80/X vssd1 vssd1 vccd1 vccd1 _1536_/X sky130_fd_sc_hd__mux2_1
XANTENNA__1372__A1 _2187_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xoutput479 hold642/X vssd1 vssd1 vccd1 vccd1 la_data_out[64] sky130_fd_sc_hd__buf_12
X_1467_ _0986_/Y hold78/X _1202_/Y hold111/X vssd1 vssd1 vccd1 vccd1 _1467_/X sky130_fd_sc_hd__a211o_1
XANTENNA__1124__A1 _2102_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_1398_ _1398_/A1 _1529_/A2 _1529_/B1 _2179_/Q hold512/X vssd1 vssd1 vccd1 vccd1 _1398_/X
+ sky130_fd_sc_hd__a221o_1
XANTENNA__1370__A _1415_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_2019_ _2033_/A vssd1 vssd1 vccd1 vccd1 _2019_/Y sky130_fd_sc_hd__inv_2
XANTENNA_fanout537_A hold79/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_45_373 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_20_207 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
Xhold160 la_data_in[47] vssd1 vssd1 vccd1 vccd1 hold93/A sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_13_281 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
Xhold171 _1474_/X vssd1 vssd1 vccd1 vccd1 _2149_/D sky130_fd_sc_hd__dlygate4sd3_1
Xhold193 la_data_in[24] vssd1 vssd1 vccd1 vccd1 hold193/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold182 hold182/A vssd1 vssd1 vccd1 vccd1 _1322_/B sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA__1115__A1 hold646/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__1280__A _1310_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_28_307 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_24_502 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_3_418 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_36_373 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_51_354 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_51_387 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_1321_ hold73/X _2204_/Q hold27/X vssd1 vssd1 vccd1 vccd1 hold74/A sky130_fd_sc_hd__mux2_1
XANTENNA__1106__A1 _2111_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_1252_ hold326/X _2227_/Q _1252_/S vssd1 vssd1 vccd1 vccd1 _1252_/X sky130_fd_sc_hd__mux2_1
X_1183_ hold625/X _1183_/A2 _1183_/B1 _1182_/X vssd1 vssd1 vccd1 vccd1 _2253_/D sky130_fd_sc_hd__a22o_1
XFILLER_0_47_605 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_19_329 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_24_73 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__1290__B1 _1529_/B1 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_55_671 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_0967_ hold35/X _0977_/B vssd1 vssd1 vccd1 vccd1 _0967_/Y sky130_fd_sc_hd__nand2_1
XFILLER_0_15_524 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_54_192 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_30_505 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__1593__B2 _2090_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xoutput276 _1753_/X vssd1 vssd1 vccd1 vccd1 data_out[111] sky130_fd_sc_hd__buf_12
Xoutput265 _1743_/X vssd1 vssd1 vccd1 vccd1 data_out[101] sky130_fd_sc_hd__buf_12
XFILLER_0_49_81 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xoutput287 _1763_/X vssd1 vssd1 vccd1 vccd1 data_out[121] sky130_fd_sc_hd__buf_12
X_1519_ _1519_/A1 _1519_/A2 _1519_/B1 _2127_/Q hold450/X vssd1 vssd1 vccd1 vccd1 _1519_/X
+ sky130_fd_sc_hd__a221o_1
Xoutput298 _1773_/X vssd1 vssd1 vccd1 vccd1 data_out[131] sky130_fd_sc_hd__buf_12
XANTENNA__1281__B1 _1527_/B1 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_52_118 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_45_181 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_21_505 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_33_365 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__1272__B1 _1519_/B1 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_1870_ _2002_/A vssd1 vssd1 vccd1 vccd1 _1870_/Y sky130_fd_sc_hd__inv_2
XFILLER_0_24_332 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XANTENNA__1575__B2 _2099_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xhold918 _1618_/X vssd1 vssd1 vccd1 vccd1 _2077_/D sky130_fd_sc_hd__dlygate4sd3_1
Xhold907 _2306_/Q vssd1 vssd1 vccd1 vccd1 hold907/X sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_12_527 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xhold929 _2100_/Q vssd1 vssd1 vccd1 vccd1 hold929/X sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA__1327__A1 _2202_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_1304_ _1310_/A hold94/X vssd1 vssd1 vccd1 vccd1 hold95/A sky130_fd_sc_hd__and2_1
XFILLER_0_19_62 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__1913__A _1913_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_2284_ _2312_/CLK _2284_/D _2023_/Y vssd1 vssd1 vccd1 vccd1 _2284_/Q sky130_fd_sc_hd__dfrtp_1
X_1235_ _1271_/A _1235_/B vssd1 vssd1 vccd1 vccd1 _1235_/X sky130_fd_sc_hd__and2_1
X_1166_ hold992/X _2081_/Q _1188_/S vssd1 vssd1 vccd1 vccd1 _1166_/X sky130_fd_sc_hd__mux2_1
X_1097_ hold572/X _1097_/A2 _1097_/B1 _1096_/X vssd1 vssd1 vccd1 vccd1 _2296_/D sky130_fd_sc_hd__a22o_1
XANTENNA__1263__B1 _1519_/B1 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_34_129 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_15_343 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_1999_ _2008_/A vssd1 vssd1 vccd1 vccd1 _1999_/Y sky130_fd_sc_hd__inv_2
XFILLER_0_42_173 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_15_376 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__1318__A1 _2205_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__1034__S _1094_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_53_405 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__1254__B1 _1503_/B1 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_46_490 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA_hold983_A _2074_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_33_140 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_34_685 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XANTENNA__1557__B2 _2108_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_21_335 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__1309__A1 _2208_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_508 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_519 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__1733__A _2171_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_1020_ hold21/X hold77/X _1192_/B hold37/X hold493/X vssd1 vssd1 vccd1 vccd1 _1020_/X
+ sky130_fd_sc_hd__o2111a_1
XANTENNA__1493__B1 _1503_/B1 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_8_307 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_29_435 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_29_446 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_1922_ _1922_/A vssd1 vssd1 vccd1 vccd1 _1922_/Y sky130_fd_sc_hd__inv_2
XFILLER_0_44_449 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_44_427 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_1853_ _1988_/A vssd1 vssd1 vccd1 vccd1 _1853_/Y sky130_fd_sc_hd__inv_2
XANTENNA__1908__A _1922_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_1784_ _2222_/Q _1798_/B vssd1 vssd1 vccd1 vccd1 _1784_/X sky130_fd_sc_hd__and2_1
XANTENNA__1548__A1 _2112_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xhold737 hold875/X vssd1 vssd1 vccd1 vccd1 hold737/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold715 hold871/X vssd1 vssd1 vccd1 vccd1 hold715/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold704 hold817/X vssd1 vssd1 vccd1 vccd1 hold704/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold726 hold855/X vssd1 vssd1 vccd1 vccd1 hold726/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold748 hold767/X vssd1 vssd1 vccd1 vccd1 hold768/A sky130_fd_sc_hd__buf_1
Xhold759 _0995_/X vssd1 vssd1 vccd1 vccd1 hold759/X sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_40_677 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_40_699 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__1643__A _2071_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_2267_ _2291_/CLK _2267_/D _2006_/Y vssd1 vssd1 vccd1 vccd1 _2267_/Q sky130_fd_sc_hd__dfrtp_1
XFILLER_0_46_93 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_1218_ input65/X _1503_/A2 _1503_/B1 _2239_/Q hold415/X vssd1 vssd1 vccd1 vccd1 _1218_/X
+ sky130_fd_sc_hd__a221o_1
XFILLER_0_27_3 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_2198_ _2219_/CLK _2198_/D _1938_/Y vssd1 vssd1 vccd1 vccd1 _2198_/Q sky130_fd_sc_hd__dfrtp_4
X_1149_ hold639/X _1183_/A2 _1183_/B1 _1148_/X vssd1 vssd1 vccd1 vccd1 _2270_/D sky130_fd_sc_hd__a22o_1
XFILLER_0_47_221 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA_fanout617_A input262/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_35_405 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_35_427 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_16_641 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_35_449 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__1539__A1 _1539_/A1 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__1539__B2 _2117_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xhold20 la_data_in[95] vssd1 vssd1 vccd1 vccd1 hold20/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold31 hold31/A vssd1 vssd1 vccd1 vccd1 hold31/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold53 hold53/A vssd1 vssd1 vccd1 vccd1 hold53/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold42 hold42/A vssd1 vssd1 vccd1 vccd1 hold42/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold64 hold64/A vssd1 vssd1 vccd1 vccd1 hold64/X sky130_fd_sc_hd__dlymetal6s2s_1
Xhold86 hold86/A vssd1 vssd1 vccd1 vccd1 hold86/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold75 la_data_in[93] vssd1 vssd1 vccd1 vccd1 hold75/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold97 hold97/A vssd1 vssd1 vccd1 vccd1 hold97/X sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_42_29 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__1227__B1 _1503_/B1 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_53_202 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_26_416 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_26_438 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_53_257 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__1728__A _2166_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_6 la_data_in[40] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_6_29 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_21_154 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_305 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_21_187 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_316 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_327 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_338 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_349 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__1463__A _2151_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_2121_ _2256_/CLK _2121_/D _1864_/Y vssd1 vssd1 vccd1 vccd1 _2121_/Q sky130_fd_sc_hd__dfrtp_4
X_2052_ _2061_/A vssd1 vssd1 vccd1 vccd1 _2052_/Y sky130_fd_sc_hd__inv_2
X_1003_ _2248_/Q _1445_/A vssd1 vssd1 vccd1 vccd1 _1003_/Y sky130_fd_sc_hd__nor2_4
XFILLER_0_16_52 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__1466__A0 _1193_/Y vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_16_63 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_16_85 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__1402__S _1435_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_9_649 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_29_243 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__1218__B1 _1503_/B1 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_17_438 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_1905_ _1913_/A vssd1 vssd1 vccd1 vccd1 _1905_/Y sky130_fd_sc_hd__inv_2
XFILLER_0_32_408 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_32_419 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_1836_ _1852_/A vssd1 vssd1 vccd1 vccd1 _1836_/Y sky130_fd_sc_hd__inv_2
Xhold501 _1266_/X vssd1 vssd1 vccd1 vccd1 hold501/X sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_4_365 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_1767_ _2205_/Q _1804_/B vssd1 vssd1 vccd1 vccd1 _1767_/X sky130_fd_sc_hd__and2_2
Xhold523 hold533/X vssd1 vssd1 vccd1 vccd1 hold523/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold545 la_data_in[88] vssd1 vssd1 vccd1 vccd1 hold545/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold534 hold538/X vssd1 vssd1 vccd1 vccd1 hold534/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold512 _1397_/Y vssd1 vssd1 vccd1 vccd1 hold512/X sky130_fd_sc_hd__buf_1
X_1698_ _2126_/Q _1715_/B vssd1 vssd1 vccd1 vccd1 _1698_/X sky130_fd_sc_hd__and2_1
Xhold556 _1194_/X vssd1 vssd1 vccd1 vccd1 _1200_/S sky130_fd_sc_hd__dlymetal6s2s_1
XFILLER_0_13_688 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xhold578 hold664/X vssd1 vssd1 vccd1 vccd1 hold578/X sky130_fd_sc_hd__dlymetal6s2s_1
Xhold567 hold678/X vssd1 vssd1 vccd1 vccd1 hold567/X sky130_fd_sc_hd__clkbuf_2
Xhold589 hold668/X vssd1 vssd1 vccd1 vccd1 hold589/X sky130_fd_sc_hd__buf_1
XANTENNA__1373__A _1415_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_861 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_850 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_894 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_883 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_872 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_2319_ _2330_/CLK _2319_/D _2058_/Y vssd1 vssd1 vccd1 vccd1 _2319_/Q sky130_fd_sc_hd__dfrtp_1
XANTENNA_fanout567_A _1003_/Y vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__1312__S _1318_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_48_585 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xcontroller_620 vssd1 vssd1 vccd1 vccd1 controller_620/HI la_data_out[2] sky130_fd_sc_hd__conb_1
Xcontroller_631 vssd1 vssd1 vccd1 vccd1 controller_631/HI la_data_out[13] sky130_fd_sc_hd__conb_1
Xcontroller_642 vssd1 vssd1 vccd1 vccd1 controller_642/HI la_data_out[24] sky130_fd_sc_hd__conb_1
XFILLER_0_50_216 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_50_205 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xcontroller_653 vssd1 vssd1 vccd1 vccd1 controller_653/HI la_data_out[117] sky130_fd_sc_hd__conb_1
XFILLER_0_43_290 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_31_430 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__1283__A _1310_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xinput110 data_in[51] vssd1 vssd1 vccd1 vccd1 _1529_/A1 sky130_fd_sc_hd__buf_1
Xinput132 data_in[71] vssd1 vssd1 vccd1 vccd1 _1489_/A1 sky130_fd_sc_hd__clkbuf_2
Xinput121 data_in[61] vssd1 vssd1 vccd1 vccd1 _1509_/A1 sky130_fd_sc_hd__clkbuf_2
Xinput143 data_in[81] vssd1 vssd1 vccd1 vccd1 _1469_/A1 sky130_fd_sc_hd__buf_1
Xinput154 data_in[91] vssd1 vssd1 vccd1 vccd1 _1419_/A1 sky130_fd_sc_hd__buf_1
Xinput176 hold519/X vssd1 vssd1 vccd1 vccd1 _1808_/C sky130_fd_sc_hd__dlymetal6s2s_1
Xinput187 hold274/X vssd1 vssd1 vccd1 vccd1 hold275/A sky130_fd_sc_hd__buf_1
Xinput165 hold52/X vssd1 vssd1 vccd1 vccd1 hold53/A sky130_fd_sc_hd__clkbuf_1
XANTENNA__1730__B _1761_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xinput198 hold189/X vssd1 vssd1 vccd1 vccd1 hold190/A sky130_fd_sc_hd__clkbuf_1
XANTENNA__1222__S _1252_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_27_703 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_1621_ _1621_/A1 _1623_/A2 _1623_/B1 _2076_/Q hold68/X vssd1 vssd1 vccd1 vccd1 _1621_/X
+ sky130_fd_sc_hd__a221o_1
XFILLER_0_34_290 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_22_474 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_22_485 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_1552_ hold192/X hold991/X _1632_/S vssd1 vssd1 vccd1 vccd1 _2110_/D sky130_fd_sc_hd__mux2_1
XANTENNA__1193__A _1810_/C vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_1483_ _1483_/A1 _1503_/A2 _1503_/B1 _2145_/Q hold443/X vssd1 vssd1 vccd1 vccd1 _1483_/X
+ sky130_fd_sc_hd__a221o_1
XTAP_124 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_146 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_135 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_157 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_179 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_168 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__1921__A _1922_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_2104_ _2168_/CLK _2104_/D _1847_/Y vssd1 vssd1 vccd1 vccd1 _2104_/Q sky130_fd_sc_hd__dfrtp_4
XANTENNA__1151__A2 _1183_/A2 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_2035_ _2065_/A vssd1 vssd1 vccd1 vccd1 _2035_/Y sky130_fd_sc_hd__inv_2
XFILLER_0_45_511 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_45_500 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_45_577 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_45_566 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_17_279 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_32_227 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_1819_ _1852_/A vssd1 vssd1 vccd1 vccd1 _1819_/Y sky130_fd_sc_hd__inv_2
XFILLER_0_13_452 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
Xhold320 _1530_/X vssd1 vssd1 vccd1 vccd1 _2121_/D sky130_fd_sc_hd__dlygate4sd3_1
Xhold342 hold376/X vssd1 vssd1 vccd1 vccd1 hold342/X sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_13_496 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xhold331 _1500_/X vssd1 vssd1 vccd1 vccd1 _2136_/D sky130_fd_sc_hd__dlygate4sd3_1
Xhold353 _1286_/X vssd1 vssd1 vccd1 vccd1 hold353/X sky130_fd_sc_hd__buf_1
Xhold386 _1490_/X vssd1 vssd1 vccd1 vccd1 _2141_/D sky130_fd_sc_hd__dlygate4sd3_1
Xhold375 hold912/X vssd1 vssd1 vccd1 vccd1 hold375/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold364 hold887/X vssd1 vssd1 vccd1 vccd1 hold364/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold397 la_data_in[71] vssd1 vssd1 vccd1 vccd1 hold397/X sky130_fd_sc_hd__dlygate4sd3_1
XTAP_691 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_680 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__1042__S _1094_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_55_308 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_36_544 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_51_558 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__1725__B _1725_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_31_293 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__1741__A _2179_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__1133__A2 _1183_/A2 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_59_614 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_0983_ hold36/X _0983_/B vssd1 vssd1 vccd1 vccd1 _0983_/Y sky130_fd_sc_hd__nor2_1
XFILLER_0_54_341 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_14_205 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_42_547 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_14_249 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
Xoutput403 _1649_/X vssd1 vssd1 vccd1 vccd1 data_out[7] sky130_fd_sc_hd__buf_12
Xoutput414 _1650_/X vssd1 vssd1 vccd1 vccd1 data_out[8] sky130_fd_sc_hd__buf_12
Xoutput425 _1651_/X vssd1 vssd1 vccd1 vccd1 data_out[9] sky130_fd_sc_hd__buf_12
X_1604_ _1603_/X _2084_/Q _1622_/S vssd1 vssd1 vccd1 vccd1 _1604_/X sky130_fd_sc_hd__mux2_1
Xoutput436 hold599/X vssd1 vssd1 vccd1 vccd1 la_data_out[109] sky130_fd_sc_hd__buf_12
XFILLER_0_10_433 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
Xoutput447 hold605/X vssd1 vssd1 vccd1 vccd1 la_data_out[32] sky130_fd_sc_hd__buf_12
Xoutput458 hold629/X vssd1 vssd1 vccd1 vccd1 la_data_out[43] sky130_fd_sc_hd__buf_12
Xoutput469 hold742/X vssd1 vssd1 vccd1 vccd1 hold743/A sky130_fd_sc_hd__buf_6
XFILLER_0_2_699 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_1535_ _1535_/A1 _1197_/D _1541_/B1 _2119_/Q hold141/X vssd1 vssd1 vccd1 vccd1 _1535_/X
+ sky130_fd_sc_hd__a221o_1
X_1466_ _1193_/Y _2152_/Q _1466_/S vssd1 vssd1 vccd1 vccd1 _1466_/X sky130_fd_sc_hd__mux2_1
X_1397_ _2249_/Q _1397_/B vssd1 vssd1 vccd1 vccd1 _1397_/Y sky130_fd_sc_hd__nor2_1
XANTENNA__1651__A _2079_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_2018_ _2033_/A vssd1 vssd1 vccd1 vccd1 _2018_/Y sky130_fd_sc_hd__inv_2
XFILLER_0_49_135 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_18_511 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_37_308 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_33_503 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_45_396 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_33_547 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_20_219 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
Xhold150 hold840/X vssd1 vssd1 vccd1 vccd1 hold47/A sky130_fd_sc_hd__dlygate4sd3_1
Xhold161 _1538_/X vssd1 vssd1 vccd1 vccd1 _2117_/D sky130_fd_sc_hd__dlygate4sd3_1
Xhold172 hold873/X vssd1 vssd1 vccd1 vccd1 hold99/A sky130_fd_sc_hd__dlygate4sd3_1
Xhold194 hold869/X vssd1 vssd1 vccd1 vccd1 hold194/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold183 _1322_/X vssd1 vssd1 vccd1 vccd1 hold183/X sky130_fd_sc_hd__buf_1
XANTENNA__1115__A2 _1183_/A2 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__1500__S _1504_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_50_29 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XANTENNA__1587__C1 hold525/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__1736__A _2174_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_1320_ input28/X _1527_/A2 _1541_/B1 _2205_/Q hold72/X vssd1 vssd1 vccd1 vccd1 hold73/A
+ sky130_fd_sc_hd__a221o_1
X_1251_ input53/X _1495_/A2 _1495_/B1 _2228_/Q hold325/X vssd1 vssd1 vccd1 vccd1 _1251_/X
+ sky130_fd_sc_hd__a221o_1
X_1182_ hold984/X _2073_/Q _1188_/S vssd1 vssd1 vccd1 vccd1 _1182_/X sky130_fd_sc_hd__mux2_1
XFILLER_0_24_85 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XANTENNA__1290__B2 _2215_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_27_363 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_6_268 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_0966_ _0978_/A _0978_/B _0971_/C _0966_/D vssd1 vssd1 vccd1 vccd1 _1455_/B sky130_fd_sc_hd__or4_2
Xclkbuf_leaf_9_wb_clk_i clkbuf_leaf_9_wb_clk_i/A vssd1 vssd1 vccd1 vccd1 _2256_/CLK
+ sky130_fd_sc_hd__clkbuf_16
XFILLER_0_42_344 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__1646__A _2074_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xoutput266 _1744_/X vssd1 vssd1 vccd1 vccd1 data_out[102] sky130_fd_sc_hd__buf_12
XFILLER_0_57_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
Xoutput277 _1754_/X vssd1 vssd1 vccd1 vccd1 data_out[112] sky130_fd_sc_hd__buf_12
Xoutput288 _1764_/X vssd1 vssd1 vccd1 vccd1 data_out[122] sky130_fd_sc_hd__buf_12
Xoutput299 _1774_/X vssd1 vssd1 vccd1 vccd1 data_out[132] sky130_fd_sc_hd__buf_12
X_1518_ _1517_/X hold945/X _1520_/S vssd1 vssd1 vccd1 vccd1 _1518_/X sky130_fd_sc_hd__mux2_1
X_1449_ _1192_/C _2160_/Q _1461_/S vssd1 vssd1 vccd1 vccd1 _1449_/X sky130_fd_sc_hd__mux2_1
XFILLER_0_38_617 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XANTENNA__1281__B2 _2218_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__1569__C1 hold244/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_33_333 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_21_517 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_45_29 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_28_105 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_29_617 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_28_116 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__1272__B2 _2221_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_37_661 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_37_694 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_52_642 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_24_344 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
Xhold919 la_data_in[6] vssd1 vssd1 vccd1 vccd1 hold62/A sky130_fd_sc_hd__dlygate4sd3_1
Xhold908 la_data_in[36] vssd1 vssd1 vccd1 vccd1 hold908/X sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_24_377 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_1303_ hold142/X _2210_/Q _1318_/S vssd1 vssd1 vccd1 vccd1 _1303_/X sky130_fd_sc_hd__mux2_1
X_2283_ _2300_/CLK _2283_/D _2022_/Y vssd1 vssd1 vccd1 vccd1 _2283_/Q sky130_fd_sc_hd__dfrtp_1
X_1234_ _1233_/X _2233_/Q _1252_/S vssd1 vssd1 vccd1 vccd1 _1234_/X sky130_fd_sc_hd__mux2_1
XANTENNA__1405__S _1435_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_1165_ hold641/X _1183_/A2 _1183_/B1 _1164_/X vssd1 vssd1 vccd1 vccd1 _2262_/D sky130_fd_sc_hd__a22o_1
XFILLER_0_35_40 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_1096_ _2208_/Q hold792/X _1112_/S vssd1 vssd1 vccd1 vccd1 _1096_/X sky130_fd_sc_hd__mux2_1
XFILLER_0_19_127 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__1263__B2 _2224_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__1263__A1 input49/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_7_511 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_51_94 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_43_631 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_1998_ _2008_/A vssd1 vssd1 vccd1 vccd1 _1998_/Y sky130_fd_sc_hd__inv_2
XFILLER_0_27_193 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_42_141 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA_fanout597_A _0952_/Y vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_11_583 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__1315__S _1318_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_clkbuf_leaf_18_wb_clk_i_A clkbuf_1_1__f_wb_clk_i/X vssd1 vssd1 vccd1 vccd1
+ sky130_fd_sc_hd__diode_2
XANTENNA__1050__S _1094_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__1254__A1 input52/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_46_480 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_18_193 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__1286__A _1310_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__1557__A2 _1623_/A2 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_hold976_A _2203_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_509 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__1225__S _1252_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__1493__A1 _1493_/A1 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_1921_ _1922_/A vssd1 vssd1 vccd1 vccd1 _1921_/Y sky130_fd_sc_hd__inv_2
XFILLER_0_29_469 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__1245__A1 input55/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_44_439 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_44_417 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_1852_ _1852_/A vssd1 vssd1 vccd1 vccd1 _1852_/Y sky130_fd_sc_hd__inv_2
XFILLER_0_25_631 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_1783_ _2221_/Q _1798_/B vssd1 vssd1 vccd1 vccd1 _1783_/X sky130_fd_sc_hd__and2_1
XFILLER_0_21_86 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_24_141 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_24_163 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xhold705 hold893/X vssd1 vssd1 vccd1 vccd1 hold705/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold727 hold845/X vssd1 vssd1 vccd1 vccd1 hold727/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold716 hold831/X vssd1 vssd1 vccd1 vccd1 hold716/X sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_40_634 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
Xhold738 hold832/X vssd1 vssd1 vccd1 vccd1 hold738/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold749 hold749/A vssd1 vssd1 vccd1 vccd1 la_data_out[122] sky130_fd_sc_hd__buf_12
XANTENNA__1924__A _1941_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__1643__B _1725_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__1181__B1 _1183_/B1 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_46_50 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_2266_ _2296_/CLK _2266_/D _2005_/Y vssd1 vssd1 vccd1 vccd1 _2266_/Q sky130_fd_sc_hd__dfrtp_1
XFILLER_0_46_83 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_2197_ _2217_/CLK _2197_/D _1937_/Y vssd1 vssd1 vccd1 vccd1 _2197_/Q sky130_fd_sc_hd__dfrtp_4
X_1217_ _1277_/A _1217_/B vssd1 vssd1 vccd1 vccd1 _1217_/X sky130_fd_sc_hd__and2_1
X_1148_ _2182_/Q _2090_/Q _1178_/S vssd1 vssd1 vccd1 vccd1 _1148_/X sky130_fd_sc_hd__mux2_1
X_1079_ hold635/X _1095_/A2 _1095_/B1 _1078_/X vssd1 vssd1 vccd1 vccd1 _2305_/D sky130_fd_sc_hd__a22o_1
XANTENNA__1236__A1 input59/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__1539__A2 _1197_/D vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_16_697 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_30_122 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_30_155 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XANTENNA__1834__A _1922_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xhold21 hold21/A vssd1 vssd1 vccd1 vccd1 hold21/X sky130_fd_sc_hd__clkbuf_2
Xhold10 la_data_in[45] vssd1 vssd1 vccd1 vccd1 hold10/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold32 hold32/A vssd1 vssd1 vccd1 vccd1 hold32/X sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA__1172__A0 _2170_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xhold65 hold65/A vssd1 vssd1 vccd1 vccd1 hold65/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold43 hold43/A vssd1 vssd1 vccd1 vccd1 hold43/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold54 hold54/A vssd1 vssd1 vccd1 vccd1 hold54/X sky130_fd_sc_hd__buf_1
Xhold87 hold87/A vssd1 vssd1 vccd1 vccd1 hold87/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold76 hold76/A vssd1 vssd1 vccd1 vccd1 hold76/X sky130_fd_sc_hd__dlymetal6s2s_1
Xhold98 hold98/A vssd1 vssd1 vccd1 vccd1 hold98/X sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA__1475__A1 _1475_/A1 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__1227__A1 input62/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_53_225 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__1728__B _1761_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_7 la_data_in[45] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__1744__A _2182_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_306 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_317 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_328 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_339 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_21_199 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XANTENNA__1163__B1 _1183_/B1 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xclkbuf_leaf_23_wb_clk_i clkbuf_1_1__f_wb_clk_i/X vssd1 vssd1 vccd1 vccd1 _2269_/CLK
+ sky130_fd_sc_hd__clkbuf_16
X_2120_ _2212_/CLK _2120_/D _1863_/Y vssd1 vssd1 vccd1 vccd1 _2120_/Q sky130_fd_sc_hd__dfrtp_4
X_2051_ _2065_/A vssd1 vssd1 vccd1 vccd1 _2051_/Y sky130_fd_sc_hd__inv_2
X_1002_ _1002_/A hold22/X vssd1 vssd1 vccd1 vccd1 _1002_/Y sky130_fd_sc_hd__nand2_1
XFILLER_0_29_222 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__1218__A1 input65/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__1919__A _1941_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_1904_ _1913_/A vssd1 vssd1 vccd1 vccd1 _1904_/Y sky130_fd_sc_hd__inv_2
XFILLER_0_29_277 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_32_85 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_1835_ _1922_/A vssd1 vssd1 vccd1 vccd1 _1835_/Y sky130_fd_sc_hd__inv_2
Xhold502 _1267_/X vssd1 vssd1 vccd1 vccd1 _2222_/D sky130_fd_sc_hd__dlygate4sd3_1
X_1766_ _2204_/Q _1766_/B vssd1 vssd1 vccd1 vccd1 _1766_/X sky130_fd_sc_hd__and2_1
Xhold513 hold517/X vssd1 vssd1 vccd1 vccd1 hold513/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold524 _1635_/B vssd1 vssd1 vccd1 vccd1 _1379_/B sky130_fd_sc_hd__dlygate4sd3_1
Xhold535 _1809_/B vssd1 vssd1 vccd1 vccd1 _1376_/B sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_4_377 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_40_431 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_1697_ _2125_/Q _1715_/B vssd1 vssd1 vccd1 vccd1 _1697_/X sky130_fd_sc_hd__and2_1
Xhold557 _1195_/X vssd1 vssd1 vccd1 vccd1 _2246_/D sky130_fd_sc_hd__dlygate4sd3_1
Xhold546 _1453_/C vssd1 vssd1 vccd1 vccd1 _0987_/D sky130_fd_sc_hd__dlygate4sd3_1
Xhold579 hold683/X vssd1 vssd1 vccd1 vccd1 hold579/X sky130_fd_sc_hd__clkbuf_2
XANTENNA__1654__A _2082_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xhold568 hold726/X vssd1 vssd1 vccd1 vccd1 hold568/X sky130_fd_sc_hd__clkbuf_2
XFILLER_0_40_464 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_40_475 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_862 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_851 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_840 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__1154__A0 _2179_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_884 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_873 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_2318_ _2328_/CLK _2318_/D _2057_/Y vssd1 vssd1 vccd1 vccd1 _2318_/Q sky130_fd_sc_hd__dfrtp_1
X_2249_ _2249_/CLK _2249_/D _1988_/Y vssd1 vssd1 vccd1 vccd1 _2249_/Q sky130_fd_sc_hd__dfrtp_2
XANTENNA__1209__A1 input69/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_36_704 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xcontroller_621 vssd1 vssd1 vccd1 vccd1 controller_621/HI la_data_out[3] sky130_fd_sc_hd__conb_1
Xcontroller_632 vssd1 vssd1 vccd1 vccd1 controller_632/HI la_data_out[14] sky130_fd_sc_hd__conb_1
XFILLER_0_35_225 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xcontroller_654 vssd1 vssd1 vccd1 vccd1 controller_654/HI la_data_out[118] sky130_fd_sc_hd__conb_1
Xcontroller_643 vssd1 vssd1 vccd1 vccd1 controller_643/HI la_data_out[25] sky130_fd_sc_hd__conb_1
XFILLER_0_23_409 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_35_258 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_31_442 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_31_475 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_9_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xinput111 data_in[52] vssd1 vssd1 vccd1 vccd1 _1527_/A1 sky130_fd_sc_hd__buf_1
Xinput100 data_in[42] vssd1 vssd1 vccd1 vccd1 _1547_/A1 sky130_fd_sc_hd__buf_1
XANTENNA__1145__B1 _1157_/B1 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xinput144 data_in[82] vssd1 vssd1 vccd1 vccd1 _1446_/A1 sky130_fd_sc_hd__buf_1
Xinput133 data_in[72] vssd1 vssd1 vccd1 vccd1 _1487_/A1 sky130_fd_sc_hd__clkbuf_2
Xinput122 data_in[62] vssd1 vssd1 vccd1 vccd1 _1507_/A1 sky130_fd_sc_hd__clkbuf_2
Xinput155 data_in[92] vssd1 vssd1 vccd1 vccd1 _1416_/A1 sky130_fd_sc_hd__buf_1
Xinput177 hold527/X vssd1 vssd1 vccd1 vccd1 _1808_/D sky130_fd_sc_hd__dlymetal6s2s_1
Xinput166 hold154/X vssd1 vssd1 vccd1 vccd1 hold155/A sky130_fd_sc_hd__clkbuf_1
Xinput199 hold181/X vssd1 vssd1 vccd1 vccd1 hold182/A sky130_fd_sc_hd__clkbuf_1
Xinput188 hold261/X vssd1 vssd1 vccd1 vccd1 hold243/A sky130_fd_sc_hd__clkbuf_1
XANTENNA__1739__A _2177_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_26_225 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__1620__A1 _2076_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_26_269 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_1620_ _1619_/X _2076_/Q _1622_/S vssd1 vssd1 vccd1 vccd1 hold82/A sky130_fd_sc_hd__mux2_1
X_1551_ input98/X _1637_/B _1635_/C _2111_/Q hold191/X vssd1 vssd1 vccd1 vccd1 _1551_/X
+ sky130_fd_sc_hd__a221o_1
X_1482_ hold516/X hold776/X _1504_/S vssd1 vssd1 vccd1 vccd1 _2145_/D sky130_fd_sc_hd__mux2_1
XANTENNA__1136__A0 _2188_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_125 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_147 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_136 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_158 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_169 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_2103_ _2194_/CLK _2103_/D _1846_/Y vssd1 vssd1 vccd1 vccd1 _2103_/Q sky130_fd_sc_hd__dfrtp_4
XFILLER_0_27_41 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_2034_ _2034_/A vssd1 vssd1 vccd1 vccd1 _2034_/Y sky130_fd_sc_hd__inv_2
XFILLER_0_43_40 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__1649__A _2077_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_9_447 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_9_436 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_45_534 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_17_225 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_45_556 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__1611__A1 input12/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__1611__B2 _2081_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_33_707 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_1818_ _1852_/A vssd1 vssd1 vccd1 vccd1 _1818_/Y sky130_fd_sc_hd__inv_2
Xhold310 hold330/X vssd1 vssd1 vccd1 vccd1 hold310/X sky130_fd_sc_hd__dlygate4sd3_1
X_1749_ _2187_/Q _1761_/B vssd1 vssd1 vccd1 vccd1 _1749_/X sky130_fd_sc_hd__and2_1
Xhold343 hold343/A vssd1 vssd1 vccd1 vccd1 _1337_/B sky130_fd_sc_hd__dlygate4sd3_1
Xhold321 la_data_in[64] vssd1 vssd1 vccd1 vccd1 hold321/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold332 la_data_in[65] vssd1 vssd1 vccd1 vccd1 hold332/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold354 _1287_/X vssd1 vssd1 vccd1 vccd1 hold354/X sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_7_73 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xhold387 la_data_in[68] vssd1 vssd1 vccd1 vccd1 hold387/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold365 la_data_in[53] vssd1 vssd1 vccd1 vccd1 hold365/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold376 hold908/X vssd1 vssd1 vccd1 vccd1 hold376/X sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_40_294 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
Xhold398 _1234_/X vssd1 vssd1 vccd1 vccd1 _2233_/D sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_0_391 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_670 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__1127__B1 _1189_/B1 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_692 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_681 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_hold422_A _1226_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_8_480 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_23_239 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__1118__A0 _2197_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_46_309 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_27_512 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_6_406 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_0982_ _1453_/D _0982_/B vssd1 vssd1 vccd1 vccd1 _1197_/B sky130_fd_sc_hd__nor2_1
XFILLER_0_27_534 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_42_537 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_42_559 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xoutput404 _1722_/X vssd1 vssd1 vccd1 vccd1 data_out[80] sky130_fd_sc_hd__buf_12
Xoutput415 _1732_/X vssd1 vssd1 vccd1 vccd1 data_out[90] sky130_fd_sc_hd__buf_12
Xoutput426 _1812_/X vssd1 vssd1 vccd1 vccd1 ki sky130_fd_sc_hd__buf_12
XFILLER_0_22_250 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_22_261 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__1408__S hold27/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_1603_ input56/X _1623_/A2 _1623_/B1 _2085_/Q hold85/X vssd1 vssd1 vccd1 vccd1 _1603_/X
+ sky130_fd_sc_hd__a221o_1
Xoutput459 hold641/X vssd1 vssd1 vccd1 vccd1 la_data_out[44] sky130_fd_sc_hd__buf_12
Xoutput437 hold587/X vssd1 vssd1 vccd1 vccd1 la_data_out[110] sky130_fd_sc_hd__buf_12
Xoutput448 hold655/X vssd1 vssd1 vccd1 vccd1 la_data_out[33] sky130_fd_sc_hd__buf_12
X_1534_ hold148/X hold930/X hold80/X vssd1 vssd1 vccd1 vccd1 _2119_/D sky130_fd_sc_hd__mux2_1
X_1465_ hold577/X _1466_/S _1057_/A2 vssd1 vssd1 vccd1 vccd1 _2153_/D sky130_fd_sc_hd__a21bo_1
X_1396_ _1395_/X hold922/X _1435_/S vssd1 vssd1 vccd1 vccd1 _2179_/D sky130_fd_sc_hd__mux2_1
XANTENNA__1651__B _1725_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_54_83 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_2017_ _2026_/A vssd1 vssd1 vccd1 vccd1 _2017_/Y sky130_fd_sc_hd__inv_2
XFILLER_0_49_169 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_18_501 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_18_523 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_18_578 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_18_589 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__1318__S _1318_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_41_581 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
Xhold162 hold178/X vssd1 vssd1 vccd1 vccd1 hold162/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold140 hold140/A vssd1 vssd1 vccd1 vccd1 _1301_/B sky130_fd_sc_hd__dlygate4sd3_1
Xhold151 la_data_in[48] vssd1 vssd1 vccd1 vccd1 hold151/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold195 hold259/X vssd1 vssd1 vccd1 vccd1 hold195/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold173 hold900/X vssd1 vssd1 vccd1 vccd1 hold52/A sky130_fd_sc_hd__dlygate4sd3_1
Xhold184 _1549_/X vssd1 vssd1 vccd1 vccd1 hold184/X sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_49_670 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_28_309 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__1289__A _1310_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_51_378 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__1228__S _1252_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__1752__A _2190_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_1250_ _1271_/A _1250_/B vssd1 vssd1 vccd1 vccd1 _1250_/X sky130_fd_sc_hd__and2_1
X_1181_ hold628/X _1183_/A2 _1183_/B1 _1180_/X vssd1 vssd1 vccd1 vccd1 _2254_/D sky130_fd_sc_hd__a22o_1
XANTENNA__1511__B1 _1519_/B1 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_19_309 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__1290__A2 _1529_/A2 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_24_97 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_0965_ _0977_/B _0977_/C _0976_/D hold35/X vssd1 vssd1 vccd1 vccd1 _0965_/X sky130_fd_sc_hd__or4b_1
XANTENNA__1927__A _1941_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_40_96 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__1646__B _1725_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xoutput267 _1745_/X vssd1 vssd1 vccd1 vccd1 data_out[103] sky130_fd_sc_hd__buf_12
XFILLER_0_49_72 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__1662__A _2090_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xoutput278 _1755_/X vssd1 vssd1 vccd1 vccd1 data_out[113] sky130_fd_sc_hd__buf_12
Xoutput289 _1765_/X vssd1 vssd1 vccd1 vccd1 data_out[123] sky130_fd_sc_hd__buf_12
X_1517_ _1517_/A1 _1529_/A2 _1529_/B1 _2128_/Q hold340/X vssd1 vssd1 vccd1 vccd1 _1517_/X
+ sky130_fd_sc_hd__a221o_1
XFILLER_0_10_264 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_1448_ _1192_/C hold78/X _1008_/Y vssd1 vssd1 vccd1 vccd1 _1461_/S sky130_fd_sc_hd__a21bo_2
XFILLER_0_4_85 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_1379_ _1394_/A _1379_/B vssd1 vssd1 vccd1 vccd1 _1379_/X sky130_fd_sc_hd__and2_1
XANTENNA_fanout542_A _1724_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_38_629 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_37_128 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__1281__A2 _1527_/A2 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__1569__B1 _1569_/B1 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_33_345 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_33_378 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_33_389 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__1048__S _1094_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_hold921_A _2102_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_29_607 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_29_629 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__1272__A2 _1519_/A2 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__1747__A _2185_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_24_301 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_37_673 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xhold909 _1339_/X vssd1 vssd1 vccd1 vccd1 _2198_/D sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_24_356 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_52_698 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_20_551 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_19_53 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_2282_ _2296_/CLK _2282_/D _2021_/Y vssd1 vssd1 vccd1 vccd1 _2282_/Q sky130_fd_sc_hd__dfrtp_1
X_1302_ input35/X _1197_/D _1527_/B1 _2211_/Q hold141/X vssd1 vssd1 vccd1 vccd1 _1302_/X
+ sky130_fd_sc_hd__a221o_1
X_1233_ input60/X _1503_/A2 _1503_/B1 _2234_/Q hold384/X vssd1 vssd1 vccd1 vccd1 _1233_/X
+ sky130_fd_sc_hd__a221o_1
X_1164_ _2174_/Q _2082_/Q _1188_/S vssd1 vssd1 vccd1 vccd1 _1164_/X sky130_fd_sc_hd__mux2_1
X_1095_ hold586/X _1095_/A2 _1095_/B1 _1094_/X vssd1 vssd1 vccd1 vccd1 _2297_/D sky130_fd_sc_hd__a22o_1
XFILLER_0_59_253 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_59_275 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__1263__A2 _1519_/A2 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_7_556 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_15_301 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_1997_ _2008_/A vssd1 vssd1 vccd1 vccd1 _1997_/Y sky130_fd_sc_hd__inv_2
XFILLER_0_27_150 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_28_662 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XANTENNA__1657__A _2085_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_15_323 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_15_334 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__1487__C1 hold348/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_38_437 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XANTENNA__1254__A2 _1503_/A2 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_19_651 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_19_673 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_34_610 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_33_153 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_34_665 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_21_337 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_33_186 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XANTENNA_clkbuf_leaf_3_wb_clk_i_A clkbuf_leaf_9_wb_clk_i/A vssd1 vssd1 vccd1 vccd1
+ sky130_fd_sc_hd__diode_2
XANTENNA_hold969_A _2095_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__1506__S _1520_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__1190__A1 _1810_/C vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__1493__A2 _1503_/A2 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_8_309 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_1920_ _1922_/A vssd1 vssd1 vccd1 vccd1 _1920_/Y sky130_fd_sc_hd__inv_2
X_1851_ _1916_/A vssd1 vssd1 vccd1 vccd1 _1851_/Y sky130_fd_sc_hd__inv_2
XFILLER_0_25_643 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_1782_ _2220_/Q _1802_/B vssd1 vssd1 vccd1 vccd1 _1782_/X sky130_fd_sc_hd__and2_1
XFILLER_0_21_98 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
Xhold728 hold867/X vssd1 vssd1 vccd1 vccd1 hold728/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold706 hold854/X vssd1 vssd1 vccd1 vccd1 hold706/X sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_24_197 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xhold717 hold818/X vssd1 vssd1 vccd1 vccd1 hold717/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold739 hold835/X vssd1 vssd1 vccd1 vccd1 hold739/X sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA__1181__A1 hold628/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_2265_ _2291_/CLK _2265_/D _2004_/Y vssd1 vssd1 vccd1 vccd1 _2265_/Q sky130_fd_sc_hd__dfrtp_1
XANTENNA__1940__A _1941_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_2196_ _2217_/CLK _2196_/D _1936_/Y vssd1 vssd1 vccd1 vccd1 _2196_/Q sky130_fd_sc_hd__dfrtp_4
XFILLER_0_46_62 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_1216_ _1215_/X _2239_/Q _1252_/S vssd1 vssd1 vccd1 vccd1 _1216_/X sky130_fd_sc_hd__mux2_1
X_1147_ hold617/X _1189_/A2 _1189_/B1 _1146_/X vssd1 vssd1 vccd1 vccd1 _2271_/D sky130_fd_sc_hd__a22o_1
X_1078_ _2217_/Q _2125_/Q _1086_/S vssd1 vssd1 vccd1 vccd1 _1078_/X sky130_fd_sc_hd__mux2_1
XFILLER_0_7_353 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_16_632 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_16_654 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_43_495 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_43_484 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_30_145 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_30_167 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_30_178 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XANTENNA__2011__A _2034_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xhold22 hold22/A vssd1 vssd1 vccd1 vccd1 hold22/X sky130_fd_sc_hd__buf_1
Xhold11 hold11/A vssd1 vssd1 vccd1 vccd1 hold11/X sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA__1172__A1 _2078_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xhold33 hold33/A vssd1 vssd1 vccd1 vccd1 hold33/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold44 hold44/A vssd1 vssd1 vccd1 vccd1 hold44/X sky130_fd_sc_hd__buf_1
Xhold55 hold55/A vssd1 vssd1 vccd1 vccd1 hold55/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold77 hold77/A vssd1 vssd1 vccd1 vccd1 hold77/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold66 hold92/X vssd1 vssd1 vccd1 vccd1 hold66/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold88 hold88/A vssd1 vssd1 vccd1 vccd1 hold88/X sky130_fd_sc_hd__clkbuf_2
Xhold99 hold99/A vssd1 vssd1 vccd1 vccd1 hold99/X sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_39_713 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__1227__A2 _1503_/A2 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_38_256 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_38_267 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_53_248 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_34_462 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA_8 la_data_in[48] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_22_613 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_21_134 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_307 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_318 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_329 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__1760__A _2198_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_2050_ _2065_/A vssd1 vssd1 vccd1 vccd1 _2050_/Y sky130_fd_sc_hd__inv_2
XFILLER_0_16_10 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_1001_ _1014_/C _0997_/X _1453_/D hold428/X vssd1 vssd1 vccd1 vccd1 _1001_/X sky130_fd_sc_hd__o2bb2a_1
XANTENNA__1218__A2 _1503_/A2 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_1903_ _1913_/A vssd1 vssd1 vccd1 vccd1 _1903_/Y sky130_fd_sc_hd__inv_2
XFILLER_0_29_289 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_44_226 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_1834_ _1922_/A vssd1 vssd1 vccd1 vccd1 _1834_/Y sky130_fd_sc_hd__inv_2
X_1765_ _2203_/Q _1766_/B vssd1 vssd1 vccd1 vccd1 _1765_/X sky130_fd_sc_hd__and2_1
XFILLER_0_40_421 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_4_389 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
Xhold514 hold514/A vssd1 vssd1 vccd1 vccd1 _1220_/B sky130_fd_sc_hd__dlygate4sd3_1
Xhold503 la_data_in[18] vssd1 vssd1 vccd1 vccd1 hold87/A sky130_fd_sc_hd__dlygate4sd3_1
Xhold536 _1376_/X vssd1 vssd1 vccd1 vccd1 hold536/X sky130_fd_sc_hd__buf_1
Xhold525 _1379_/X vssd1 vssd1 vccd1 vccd1 hold525/X sky130_fd_sc_hd__dlymetal6s2s_1
X_1696_ _2124_/Q _1715_/B vssd1 vssd1 vccd1 vccd1 _1696_/X sky130_fd_sc_hd__and2_1
Xhold547 _0983_/B vssd1 vssd1 vccd1 vccd1 _0982_/B sky130_fd_sc_hd__dlygate4sd3_1
Xhold558 la_data_in[84] vssd1 vssd1 vccd1 vccd1 hold558/X sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA__1654__B _1725_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xhold569 _1133_/X vssd1 vssd1 vccd1 vccd1 _2278_/D sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_0_573 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_852 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_57_50 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_841 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_830 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__1154__A1 _2087_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_885 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_874 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_863 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_2317_ _2328_/CLK _2317_/D _2056_/Y vssd1 vssd1 vccd1 vccd1 _2317_/Q sky130_fd_sc_hd__dfrtp_1
XANTENNA__1670__A _2098_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_2248_ _2249_/CLK _2248_/D _1987_/Y vssd1 vssd1 vccd1 vccd1 _2248_/Q sky130_fd_sc_hd__dfrtp_4
XFILLER_0_32_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_2179_ _2194_/CLK _2179_/D _1919_/Y vssd1 vssd1 vccd1 vccd1 _2179_/Q sky130_fd_sc_hd__dfrtp_4
Xcontroller_622 vssd1 vssd1 vccd1 vccd1 controller_622/HI la_data_out[4] sky130_fd_sc_hd__conb_1
Xcontroller_633 vssd1 vssd1 vccd1 vccd1 controller_633/HI la_data_out[15] sky130_fd_sc_hd__conb_1
Xcontroller_644 vssd1 vssd1 vccd1 vccd1 controller_644/HI la_data_out[26] sky130_fd_sc_hd__conb_1
Xcontroller_655 vssd1 vssd1 vccd1 vccd1 controller_655/HI la_data_out[119] sky130_fd_sc_hd__conb_1
XFILLER_0_31_410 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_31_487 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_12_690 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__1056__S _1094_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xinput101 data_in[43] vssd1 vssd1 vccd1 vccd1 _1545_/A1 sky130_fd_sc_hd__buf_1
Xinput134 data_in[73] vssd1 vssd1 vccd1 vccd1 _1485_/A1 sky130_fd_sc_hd__buf_2
Xinput145 data_in[83] vssd1 vssd1 vccd1 vccd1 _1443_/A1 sky130_fd_sc_hd__buf_1
Xinput112 data_in[53] vssd1 vssd1 vccd1 vccd1 _1525_/A1 sky130_fd_sc_hd__buf_1
Xinput123 data_in[63] vssd1 vssd1 vccd1 vccd1 _1505_/A1 sky130_fd_sc_hd__clkbuf_2
Xinput156 data_in[93] vssd1 vssd1 vccd1 vccd1 _1413_/A1 sky130_fd_sc_hd__buf_1
Xinput178 hold523/X vssd1 vssd1 vccd1 vccd1 _1635_/B sky130_fd_sc_hd__dlymetal6s2s_1
Xinput167 hold201/X vssd1 vssd1 vccd1 vccd1 hold202/A sky130_fd_sc_hd__clkbuf_1
Xinput189 hold404/X vssd1 vssd1 vccd1 vccd1 _1806_/B sky130_fd_sc_hd__buf_1
XFILLER_0_39_554 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__1739__B _1761_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__1081__B1 _1095_/B1 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_41_229 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_34_270 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__1755__A _2193_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_1550_ hold184/X hold989/X _1632_/S vssd1 vssd1 vccd1 vccd1 _2111_/D sky130_fd_sc_hd__mux2_1
XFILLER_0_22_421 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_34_281 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_1481_ _1481_/A1 _1503_/A2 _1503_/B1 _2146_/Q hold515/X vssd1 vssd1 vccd1 vccd1 _1481_/X
+ sky130_fd_sc_hd__a221o_1
XANTENNA__1136__A1 _2096_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_148 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_126 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_137 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_159 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_2102_ _2182_/CLK _2102_/D _1845_/Y vssd1 vssd1 vccd1 vccd1 _2102_/Q sky130_fd_sc_hd__dfrtp_4
XFILLER_0_27_75 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_2033_ _2033_/A vssd1 vssd1 vccd1 vccd1 _2033_/Y sky130_fd_sc_hd__inv_2
XFILLER_0_9_404 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_43_96 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__1072__A0 _2220_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_17_237 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_17_259 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__1611__A2 _1637_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_25_270 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_1817_ _1852_/A vssd1 vssd1 vccd1 vccd1 _1817_/Y sky130_fd_sc_hd__inv_2
XANTENNA__1665__A _2093_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xhold300 _1478_/X vssd1 vssd1 vccd1 vccd1 _2147_/D sky130_fd_sc_hd__dlygate4sd3_1
Xhold311 hold311/A vssd1 vssd1 vccd1 vccd1 _1247_/B sky130_fd_sc_hd__dlygate4sd3_1
X_1748_ _2186_/Q _1761_/B vssd1 vssd1 vccd1 vccd1 _1748_/X sky130_fd_sc_hd__and2_1
Xhold344 _1337_/X vssd1 vssd1 vccd1 vccd1 hold344/X sky130_fd_sc_hd__buf_1
Xhold333 _1502_/X vssd1 vssd1 vccd1 vccd1 _2135_/D sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA__1375__A1 _2186_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_40_251 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xhold322 _1504_/X vssd1 vssd1 vccd1 vccd1 _2134_/D sky130_fd_sc_hd__dlygate4sd3_1
Xhold366 _1526_/X vssd1 vssd1 vccd1 vccd1 _2123_/D sky130_fd_sc_hd__dlygate4sd3_1
Xhold355 _1288_/X vssd1 vssd1 vccd1 vccd1 _2215_/D sky130_fd_sc_hd__dlygate4sd3_1
X_1679_ _2107_/Q _1680_/B vssd1 vssd1 vccd1 vccd1 _1679_/X sky130_fd_sc_hd__and2_1
Xhold377 hold395/X vssd1 vssd1 vccd1 vccd1 hold377/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold399 hold439/X vssd1 vssd1 vccd1 vccd1 hold399/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold388 _1496_/X vssd1 vssd1 vccd1 vccd1 _2138_/D sky130_fd_sc_hd__dlygate4sd3_1
XTAP_660 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__1127__B2 _1126_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_693 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_682 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_671 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_fanout572_A _1201_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_48_340 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA_hold415_A _1217_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_8_470 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__1063__B1 _1097_/B1 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_hold951_A _2074_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__1118__A1 _2105_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__1514__S _1520_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_13_22 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_0981_ _1453_/B _0987_/D _1453_/A _0987_/B vssd1 vssd1 vccd1 vccd1 _0983_/B sky130_fd_sc_hd__or4bb_2
XFILLER_0_54_332 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_6_418 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_15_708 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_54_387 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_54_376 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_54_365 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_14_229 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_1602_ _1601_/X hold942/X _1622_/S vssd1 vssd1 vccd1 vccd1 _1602_/X sky130_fd_sc_hd__mux2_1
Xoutput416 _1733_/X vssd1 vssd1 vccd1 vccd1 data_out[91] sky130_fd_sc_hd__buf_12
Xoutput405 _1723_/X vssd1 vssd1 vccd1 vccd1 data_out[81] sky130_fd_sc_hd__buf_12
Xoutput438 hold588/X vssd1 vssd1 vccd1 vccd1 la_data_out[111] sky130_fd_sc_hd__buf_12
Xoutput427 hold591/X vssd1 vssd1 vccd1 vccd1 la_data_out[100] sky130_fd_sc_hd__buf_12
Xoutput449 hold603/X vssd1 vssd1 vccd1 vccd1 la_data_out[34] sky130_fd_sc_hd__buf_12
X_1533_ _1533_/A1 _1533_/A2 _1533_/B1 _2120_/Q hold147/X vssd1 vssd1 vccd1 vccd1 _1533_/X
+ sky130_fd_sc_hd__a221o_1
X_1464_ _1463_/X _2154_/Q _1464_/S vssd1 vssd1 vccd1 vccd1 _1464_/X sky130_fd_sc_hd__mux2_1
XFILLER_0_38_41 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_1395_ _1395_/A1 _1569_/A2 _1569_/B1 _2180_/Q _1394_/X vssd1 vssd1 vccd1 vccd1 _1395_/X
+ sky130_fd_sc_hd__a221o_1
XFILLER_0_54_73 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_2016_ _2034_/A vssd1 vssd1 vccd1 vccd1 _2016_/Y sky130_fd_sc_hd__inv_2
XANTENNA__1293__B1 _1529_/B1 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__1045__B1 _1095_/B1 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_18_546 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_18_568 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xhold130 hold138/X vssd1 vssd1 vccd1 vccd1 hold130/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold141 _1301_/X vssd1 vssd1 vccd1 vccd1 hold141/X sky130_fd_sc_hd__buf_1
Xhold152 _1536_/X vssd1 vssd1 vccd1 vccd1 _2118_/D sky130_fd_sc_hd__dlygate4sd3_1
Xhold174 hold213/X vssd1 vssd1 vccd1 vccd1 hold174/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold163 hold163/A vssd1 vssd1 vccd1 vccd1 _1295_/B sky130_fd_sc_hd__dlygate4sd3_1
Xhold185 hold205/X vssd1 vssd1 vccd1 vccd1 hold185/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold196 hold196/A vssd1 vssd1 vccd1 vccd1 _1313_/B sky130_fd_sc_hd__dlygate4sd3_1
Xfanout610 _2026_/A vssd1 vssd1 vccd1 vccd1 _2002_/A sky130_fd_sc_hd__buf_8
XANTENNA__1520__A1 _2126_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_490 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__1284__B1 _1529_/B1 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_48_181 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__1587__B2 _2093_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_24_505 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_51_335 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_51_357 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__1339__A1 _2198_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__1752__B _1761_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_1180_ hold979/X hold983/X _1188_/S vssd1 vssd1 vccd1 vccd1 _1180_/X sky130_fd_sc_hd__mux2_1
XANTENNA__1511__A1 _1511_/A1 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_46_107 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__1275__B1 _1529_/B1 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_24_76 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_54_173 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_0964_ _1453_/A _0987_/B _1453_/B _0987_/D vssd1 vssd1 vccd1 vccd1 _0973_/C sky130_fd_sc_hd__or4_1
XFILLER_0_15_505 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_15_527 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_40_75 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_30_508 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
Xoutput268 _1746_/X vssd1 vssd1 vccd1 vccd1 data_out[104] sky130_fd_sc_hd__buf_12
XFILLER_0_49_40 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_1516_ hold471/X _2128_/Q _1520_/S vssd1 vssd1 vccd1 vccd1 _1516_/X sky130_fd_sc_hd__mux2_1
XANTENNA__1943__A _1949_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xoutput279 _1756_/X vssd1 vssd1 vccd1 vccd1 data_out[114] sky130_fd_sc_hd__buf_12
XFILLER_0_49_84 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_1447_ _1446_/X _2162_/Q hold27/X vssd1 vssd1 vccd1 vccd1 _1447_/X sky130_fd_sc_hd__mux2_1
X_1378_ hold537/X hold986/X hold26/X vssd1 vssd1 vccd1 vccd1 _2185_/D sky130_fd_sc_hd__mux2_1
XANTENNA__1266__B1 _1519_/B1 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_18_343 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__1569__B2 _2102_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_18_365 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA_hold113_A hold79/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_33_357 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__1257__B1 _1519_/B1 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__1009__B1 _1810_/C vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_51_121 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_36_195 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_12_508 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xclkbuf_leaf_17_wb_clk_i clkbuf_1_1__f_wb_clk_i/X vssd1 vssd1 vccd1 vccd1 _2315_/CLK
+ sky130_fd_sc_hd__clkbuf_16
XFILLER_0_32_390 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__1763__A _2201_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_2281_ _2291_/CLK _2281_/D _2020_/Y vssd1 vssd1 vccd1 vccd1 _2281_/Q sky130_fd_sc_hd__dfrtp_1
X_1301_ _1310_/A _1301_/B vssd1 vssd1 vccd1 vccd1 _1301_/X sky130_fd_sc_hd__and2_1
XFILLER_0_19_65 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_1232_ _1271_/A _1232_/B vssd1 vssd1 vccd1 vccd1 _1232_/X sky130_fd_sc_hd__and2_1
X_1163_ hold640/X _1183_/A2 _1183_/B1 _1162_/X vssd1 vssd1 vccd1 vccd1 _2263_/D sky130_fd_sc_hd__a22o_1
X_1094_ _2209_/Q _2117_/Q _1094_/S vssd1 vssd1 vccd1 vccd1 _1094_/X sky130_fd_sc_hd__mux2_1
XFILLER_0_47_449 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_51_74 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_1996_ _2008_/A vssd1 vssd1 vccd1 vccd1 _1996_/Y sky130_fd_sc_hd__inv_2
XFILLER_0_28_674 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_43_622 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_27_173 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_28_696 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_15_379 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_42_176 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__1673__A _2101_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__1487__B1 _1503_/B1 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__2009__A _2034_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_38_405 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_38_449 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_46_471 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_19_685 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_33_121 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_33_165 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_34_699 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_33_198 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__1522__S hold80/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_29_427 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__1758__A _2196_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_1850_ _1916_/A vssd1 vssd1 vccd1 vccd1 _1850_/Y sky130_fd_sc_hd__inv_2
XFILLER_0_24_121 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_1781_ _2219_/Q _1798_/B vssd1 vssd1 vccd1 vccd1 _1781_/X sky130_fd_sc_hd__and2_1
XFILLER_0_4_549 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_25_655 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
Xhold718 hold872/X vssd1 vssd1 vccd1 vccd1 hold718/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold707 hold896/X vssd1 vssd1 vccd1 vccd1 hold707/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold729 hold816/X vssd1 vssd1 vccd1 vccd1 hold729/X sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_40_658 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__1181__A2 _1183_/A2 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_2264_ _2291_/CLK _2264_/D _2003_/Y vssd1 vssd1 vccd1 vccd1 _2264_/Q sky130_fd_sc_hd__dfrtp_1
X_2195_ _2217_/CLK _2195_/D _1935_/Y vssd1 vssd1 vccd1 vccd1 _2195_/Q sky130_fd_sc_hd__dfrtp_4
X_1215_ input66/X _1495_/A2 _1495_/B1 _2240_/Q hold298/X vssd1 vssd1 vccd1 vccd1 _1215_/X
+ sky130_fd_sc_hd__a221o_1
XANTENNA__1432__S _1435_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_1146_ _2183_/Q _2091_/Q _1178_/S vssd1 vssd1 vccd1 vccd1 _1146_/X sky130_fd_sc_hd__mux2_1
X_1077_ hold632/X _1095_/A2 _1095_/B1 _1076_/X vssd1 vssd1 vccd1 vccd1 _2306_/D sky130_fd_sc_hd__a22o_1
XANTENNA__1668__A _2096_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_47_246 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_1979_ _1979_/A vssd1 vssd1 vccd1 vccd1 _1979_/Y sky130_fd_sc_hd__inv_2
XFILLER_0_7_387 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_43_474 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xhold23 hold23/A vssd1 vssd1 vccd1 vccd1 hold23/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold12 hold12/A vssd1 vssd1 vccd1 vccd1 hold12/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold34 la_data_in[82] vssd1 vssd1 vccd1 vccd1 hold34/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold45 hold45/A vssd1 vssd1 vccd1 vccd1 hold45/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold56 hold56/A vssd1 vssd1 vccd1 vccd1 hold56/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold78 hold78/A vssd1 vssd1 vccd1 vccd1 hold78/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold89 hold89/A vssd1 vssd1 vccd1 vccd1 hold89/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold67 hold67/A vssd1 vssd1 vccd1 vccd1 hold67/X sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_38_213 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA_hold981_A _2092_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_9 la_data_in[52] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_22_625 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_21_124 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_21_157 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_308 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_319 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__1163__A2 _1183_/A2 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__1760__B _1761_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__1252__S _1252_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_1000_ hold22/X vssd1 vssd1 vccd1 vccd1 hold23/A sky130_fd_sc_hd__inv_2
X_1902_ _1913_/A vssd1 vssd1 vccd1 vccd1 _1902_/Y sky130_fd_sc_hd__inv_2
XFILLER_0_32_32 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__1623__B1 _1623_/B1 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_1833_ _1922_/A vssd1 vssd1 vccd1 vccd1 _1833_/Y sky130_fd_sc_hd__inv_2
X_1764_ _2202_/Q _1766_/B vssd1 vssd1 vccd1 vccd1 _1764_/X sky130_fd_sc_hd__and2_2
Xhold526 _1587_/X vssd1 vssd1 vccd1 vccd1 hold526/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold504 hold87/X vssd1 vssd1 vccd1 vccd1 hold504/X sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_25_496 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xhold515 _1220_/X vssd1 vssd1 vccd1 vccd1 hold515/X sky130_fd_sc_hd__dlymetal6s2s_1
X_1695_ _2123_/Q _1715_/B vssd1 vssd1 vccd1 vccd1 _1695_/X sky130_fd_sc_hd__and2_1
Xhold548 _1197_/B vssd1 vssd1 vccd1 vccd1 hold548/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold559 _0977_/D vssd1 vssd1 vccd1 vccd1 _0976_/D sky130_fd_sc_hd__dlygate4sd3_1
Xhold537 _1377_/X vssd1 vssd1 vccd1 vccd1 hold537/X sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_40_477 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_853 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_842 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_831 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_820 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_886 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_875 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_864 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_2316_ _2330_/CLK _2316_/D _2055_/Y vssd1 vssd1 vccd1 vccd1 _2316_/Q sky130_fd_sc_hd__dfrtp_1
X_2247_ _2249_/CLK _2247_/D _1986_/Y vssd1 vssd1 vccd1 vccd1 _2247_/Q sky130_fd_sc_hd__dfrtp_2
XANTENNA__1162__S _1188_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_25_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_2178_ _2219_/CLK _2178_/D _1918_/Y vssd1 vssd1 vccd1 vccd1 _2178_/Q sky130_fd_sc_hd__dfrtp_4
X_1129_ _2280_/Q _1189_/A2 _1189_/B1 _1128_/X vssd1 vssd1 vccd1 vccd1 _1129_/X sky130_fd_sc_hd__a22o_1
Xcontroller_623 vssd1 vssd1 vccd1 vccd1 controller_623/HI la_data_out[5] sky130_fd_sc_hd__conb_1
XANTENNA_fanout615_A input262/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__1090__A1 _2119_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xcontroller_645 vssd1 vssd1 vccd1 vccd1 controller_645/HI la_data_out[27] sky130_fd_sc_hd__conb_1
Xcontroller_634 vssd1 vssd1 vccd1 vccd1 controller_634/HI la_data_out[16] sky130_fd_sc_hd__conb_1
Xcontroller_656 vssd1 vssd1 vccd1 vccd1 controller_656/HI la_data_out[120] sky130_fd_sc_hd__conb_1
XFILLER_0_50_208 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_43_260 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__2022__A _2026_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xinput102 data_in[44] vssd1 vssd1 vccd1 vccd1 _1543_/A1 sky130_fd_sc_hd__buf_1
XANTENNA__1145__A2 _1157_/A2 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__1861__A _1941_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xinput124 data_in[64] vssd1 vssd1 vccd1 vccd1 _1503_/A1 sky130_fd_sc_hd__clkbuf_2
Xinput113 data_in[54] vssd1 vssd1 vccd1 vccd1 _1523_/A1 sky130_fd_sc_hd__buf_1
Xinput135 data_in[74] vssd1 vssd1 vccd1 vccd1 _1483_/A1 sky130_fd_sc_hd__buf_2
Xinput157 data_in[94] vssd1 vssd1 vccd1 vccd1 _1410_/A1 sky130_fd_sc_hd__buf_1
Xinput146 data_in[84] vssd1 vssd1 vccd1 vccd1 _1440_/A1 sky130_fd_sc_hd__buf_1
Xinput168 hold217/X vssd1 vssd1 vccd1 vccd1 hold218/A sky130_fd_sc_hd__buf_1
Xinput179 hold534/X vssd1 vssd1 vccd1 vccd1 _1809_/B sky130_fd_sc_hd__dlymetal6s2s_1
XANTENNA_clkbuf_1_1__f_wb_clk_i_A clkbuf_0_wb_clk_i/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__1605__B1 _1623_/B1 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__1081__B2 _1080_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_22_433 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_22_466 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_22_477 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_1480_ _1479_/X _2146_/Q _1504_/S vssd1 vssd1 vccd1 vccd1 _1480_/X sky130_fd_sc_hd__mux2_1
XFILLER_0_22_488 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_127 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_138 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__1771__A _2209_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_149 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_2101_ _2182_/CLK _2101_/D _1844_/Y vssd1 vssd1 vccd1 vccd1 _2101_/Q sky130_fd_sc_hd__dfrtp_4
X_2032_ _2033_/A vssd1 vssd1 vccd1 vccd1 _2032_/Y sky130_fd_sc_hd__inv_2
XFILLER_0_27_87 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_43_53 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_45_503 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_45_525 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_45_569 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__1946__A _1949_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_1816_ _1988_/A vssd1 vssd1 vccd1 vccd1 _1816_/Y sky130_fd_sc_hd__inv_2
Xhold301 hold915/X vssd1 vssd1 vccd1 vccd1 hold301/X sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_4_154 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_1747_ _2185_/Q _1756_/B vssd1 vssd1 vccd1 vccd1 _1747_/X sky130_fd_sc_hd__and2_1
Xhold334 hold364/X vssd1 vssd1 vccd1 vccd1 hold334/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold323 hold332/X vssd1 vssd1 vccd1 vccd1 hold323/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold312 _1247_/X vssd1 vssd1 vccd1 vccd1 hold312/X sky130_fd_sc_hd__buf_1
X_1678_ _2106_/Q _1680_/B vssd1 vssd1 vccd1 vccd1 _1678_/X sky130_fd_sc_hd__and2_1
Xhold345 _1559_/X vssd1 vssd1 vccd1 vccd1 hold345/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold378 hold378/A vssd1 vssd1 vccd1 vccd1 _1244_/B sky130_fd_sc_hd__dlygate4sd3_1
Xhold356 la_data_in[57] vssd1 vssd1 vccd1 vccd1 hold356/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold367 hold375/X vssd1 vssd1 vccd1 vccd1 hold367/X sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_13_499 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
Xhold389 hold394/X vssd1 vssd1 vccd1 vccd1 hold389/X sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA__1681__A _2109_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_661 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_650 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__1127__A2 _1189_/A2 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_694 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_683 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_672 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_fanout565_A _1529_/A2 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__2017__A _2026_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_36_547 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XANTENNA__1856__A _1913_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_16_271 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
Xhold890 _1604_/X vssd1 vssd1 vccd1 vccd1 _2084_/D sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA_hold944_A _2192_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_59_617 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_58_149 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_27_503 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_0980_ _1453_/B _0980_/B hold540/A vssd1 vssd1 vccd1 vccd1 _0980_/X sky130_fd_sc_hd__or3b_1
XANTENNA_output484_A hold646/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_27_558 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_27_569 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XANTENNA__1766__A _2204_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_1601_ input67/X _1623_/A2 _1623_/B1 _2086_/Q hold132/X vssd1 vssd1 vccd1 vccd1 _1601_/X
+ sky130_fd_sc_hd__a221o_1
Xoutput406 _1724_/X vssd1 vssd1 vccd1 vccd1 data_out[82] sky130_fd_sc_hd__buf_12
Xoutput417 _1734_/X vssd1 vssd1 vccd1 vccd1 data_out[92] sky130_fd_sc_hd__buf_12
Xoutput439 hold583/X vssd1 vssd1 vccd1 vccd1 la_data_out[112] sky130_fd_sc_hd__buf_12
Xoutput428 hold592/X vssd1 vssd1 vccd1 vccd1 la_data_out[101] sky130_fd_sc_hd__buf_12
X_1532_ _1531_/X _2120_/Q hold80/X vssd1 vssd1 vccd1 vccd1 _1532_/X sky130_fd_sc_hd__mux2_1
X_1463_ _2151_/Q _1463_/B vssd1 vssd1 vccd1 vccd1 _1463_/X sky130_fd_sc_hd__and2_1
XFILLER_0_22_296 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_1394_ _1394_/A _1394_/B vssd1 vssd1 vccd1 vccd1 _1394_/X sky130_fd_sc_hd__and2_1
XFILLER_0_38_75 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_54_41 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_2015_ _2033_/A vssd1 vssd1 vccd1 vccd1 _2015_/Y sky130_fd_sc_hd__inv_2
XFILLER_0_54_85 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_49_116 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__1293__B2 _2214_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__1676__A _2104_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_45_399 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_26_580 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_41_561 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_41_594 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xhold120 _1810_/A vssd1 vssd1 vccd1 vccd1 _1394_/B sky130_fd_sc_hd__dlygate4sd3_1
Xhold131 hold131/A vssd1 vssd1 vccd1 vccd1 _1400_/B sky130_fd_sc_hd__dlygate4sd3_1
Xhold153 la_data_in[34] vssd1 vssd1 vccd1 vccd1 hold153/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold142 _1302_/X vssd1 vssd1 vccd1 vccd1 hold142/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold186 hold186/A vssd1 vssd1 vccd1 vccd1 _1421_/B sky130_fd_sc_hd__dlygate4sd3_1
Xhold175 hold175/A vssd1 vssd1 vccd1 vccd1 _1436_/B sky130_fd_sc_hd__dlygate4sd3_1
Xhold164 _1295_/X vssd1 vssd1 vccd1 vccd1 hold164/X sky130_fd_sc_hd__buf_1
Xfanout611 input262/X vssd1 vssd1 vccd1 vccd1 _2026_/A sky130_fd_sc_hd__buf_4
Xhold197 _1313_/X vssd1 vssd1 vccd1 vccd1 hold197/X sky130_fd_sc_hd__buf_1
Xfanout600 _1922_/A vssd1 vssd1 vccd1 vccd1 _1852_/A sky130_fd_sc_hd__buf_8
XTAP_480 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_491 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__1284__B2 _2217_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_48_193 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_36_399 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_20_701 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XANTENNA__1511__A2 _1519_/A2 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_59_447 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__1275__B2 _2220_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_54_130 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_54_152 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_54_141 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_6_227 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_0963_ _0978_/A _0978_/B vssd1 vssd1 vccd1 vccd1 _0973_/B sky130_fd_sc_hd__or2_2
XFILLER_0_27_355 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_40_54 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_42_347 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_42_358 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_23_561 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_1515_ _1515_/A1 _1519_/A2 _1519_/B1 _2129_/Q hold470/X vssd1 vssd1 vccd1 vccd1 _1515_/X
+ sky130_fd_sc_hd__a221o_1
XFILLER_0_10_233 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_10_222 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xoutput269 _1747_/X vssd1 vssd1 vccd1 vccd1 data_out[105] sky130_fd_sc_hd__buf_12
XANTENNA__1435__S _1435_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_1446_ _1446_/A1 _1198_/A _1545_/B1 _2163_/Q hold49/X vssd1 vssd1 vccd1 vccd1 _1446_/X
+ sky130_fd_sc_hd__a221o_1
X_1377_ input7/X _1533_/A2 _1533_/B1 _2186_/Q hold536/X vssd1 vssd1 vccd1 vccd1 _1377_/X
+ sky130_fd_sc_hd__a221o_1
XANTENNA__1170__S _1188_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__1266__B2 _2223_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout528_A _1157_/A2 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__1569__A2 _1569_/A2 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_45_163 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_18_399 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_5_293 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__1345__S _1435_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__1257__A1 input51/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_36_163 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_37_697 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_20_531 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__1255__S hold26/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_19_11 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_2280_ _2291_/CLK _2280_/D _2019_/Y vssd1 vssd1 vccd1 vccd1 _2280_/Q sky130_fd_sc_hd__dfrtp_1
X_1300_ _1299_/X _2211_/Q _1318_/S vssd1 vssd1 vccd1 vccd1 _1300_/X sky130_fd_sc_hd__mux2_1
X_1231_ _1230_/X _2234_/Q _1252_/S vssd1 vssd1 vccd1 vccd1 _1231_/X sky130_fd_sc_hd__mux2_1
X_1162_ _2175_/Q _2083_/Q _1188_/S vssd1 vssd1 vccd1 vccd1 _1162_/X sky130_fd_sc_hd__mux2_1
X_1093_ hold579/X _1097_/A2 _1097_/B1 _1092_/X vssd1 vssd1 vccd1 vccd1 _2298_/D sky130_fd_sc_hd__a22o_1
XANTENNA__1248__A1 input54/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_47_439 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_51_86 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_43_601 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_1995_ _2002_/A vssd1 vssd1 vccd1 vccd1 _1995_/Y sky130_fd_sc_hd__inv_2
XFILLER_0_43_645 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_43_634 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_27_196 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_15_369 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__1420__A1 _2171_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__1184__A0 _2164_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_55_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_1429_ hold65/X _2168_/Q _1435_/S vssd1 vssd1 vccd1 vccd1 _1429_/X sky130_fd_sc_hd__mux2_1
XANTENNA__1487__A1 _1487_/A1 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__1239__A1 input58/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_38_417 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_19_697 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_33_111 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__2025__A _2026_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__1411__A1 _2174_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_33_133 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_21_317 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_14_391 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XANTENNA__1175__B1 _1189_/B1 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__1478__A1 _2147_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_29_406 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__1758__B _1761_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_37_461 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_1780_ _2218_/Q _1798_/B vssd1 vssd1 vccd1 vccd1 _1780_/X sky130_fd_sc_hd__and2_1
XFILLER_0_21_23 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_25_667 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
Xhold719 hold880/X vssd1 vssd1 vccd1 vccd1 hold719/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold708 hold865/X vssd1 vssd1 vccd1 vccd1 hold708/X sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA__1774__A _2212_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_0_712 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_20_394 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_2263_ _2296_/CLK _2263_/D _2002_/Y vssd1 vssd1 vccd1 vccd1 _2263_/Q sky130_fd_sc_hd__dfrtp_1
X_2194_ _2194_/CLK _2194_/D _1934_/Y vssd1 vssd1 vccd1 vccd1 _2194_/Q sky130_fd_sc_hd__dfrtp_4
X_1214_ _1277_/A _1214_/B vssd1 vssd1 vccd1 vccd1 _1214_/X sky130_fd_sc_hd__and2_1
XANTENNA__1469__A1 _1469_/A1 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_46_97 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_1145_ _2272_/Q _1157_/A2 _1157_/B1 _1144_/X vssd1 vssd1 vccd1 vccd1 _1145_/X sky130_fd_sc_hd__a22o_1
X_1076_ _2218_/Q _2126_/Q _1086_/S vssd1 vssd1 vccd1 vccd1 _1076_/X sky130_fd_sc_hd__mux2_2
XANTENNA__1949__A _1949_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_7_333 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_28_450 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_28_461 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_35_409 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_1978_ _2039_/A vssd1 vssd1 vccd1 vccd1 _1978_/Y sky130_fd_sc_hd__inv_2
XFILLER_0_16_645 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__1684__A _2112_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_31_615 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_15_199 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_30_125 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__1157__B1 _1157_/B1 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_11_383 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA_fanout595_A _1310_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xhold13 hold13/A vssd1 vssd1 vccd1 vccd1 hold13/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold24 hold24/A vssd1 vssd1 vccd1 vccd1 hold24/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold35 hold35/A vssd1 vssd1 vccd1 vccd1 hold35/X sky130_fd_sc_hd__dlymetal6s2s_1
Xhold46 hold46/A vssd1 vssd1 vccd1 vccd1 hold46/X sky130_fd_sc_hd__dlygate4sd3_1
Xclkbuf_leaf_2_wb_clk_i clkbuf_leaf_9_wb_clk_i/A vssd1 vssd1 vccd1 vccd1 _2177_/CLK
+ sky130_fd_sc_hd__clkbuf_16
Xhold57 hold57/A vssd1 vssd1 vccd1 vccd1 hold57/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold79 hold79/A vssd1 vssd1 vccd1 vccd1 hold79/X sky130_fd_sc_hd__clkbuf_2
Xhold68 hold68/A vssd1 vssd1 vccd1 vccd1 hold68/X sky130_fd_sc_hd__buf_1
XANTENNA__1859__A _1949_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_53_206 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__1632__A1 _2070_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_53_239 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_53_228 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_21_103 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_22_604 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_34_475 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_22_637 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA_hold974_A _2219_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__1148__A0 _2182_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_21_147 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_21_169 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_309 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__1320__B1 _1541_/B1 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_57_501 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__1769__A _2207_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_1901_ _1949_/A vssd1 vssd1 vccd1 vccd1 _1901_/Y sky130_fd_sc_hd__inv_2
XANTENNA__1623__B2 _2075_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_1832_ _1922_/A vssd1 vssd1 vccd1 vccd1 _1832_/Y sky130_fd_sc_hd__inv_2
XFILLER_0_44_206 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XANTENNA_clkbuf_leaf_17_wb_clk_i_A clkbuf_1_1__f_wb_clk_i/X vssd1 vssd1 vccd1 vccd1
+ sky130_fd_sc_hd__diode_2
XFILLER_0_25_486 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_1763_ _2201_/Q _1766_/B vssd1 vssd1 vccd1 vccd1 _1763_/X sky130_fd_sc_hd__and2_1
X_1694_ _2122_/Q _1715_/B vssd1 vssd1 vccd1 vccd1 _1694_/X sky130_fd_sc_hd__and2_1
Xhold505 la_data_in[60] vssd1 vssd1 vccd1 vccd1 hold505/X sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_13_637 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xhold527 hold532/X vssd1 vssd1 vccd1 vccd1 hold527/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold516 _1481_/X vssd1 vssd1 vccd1 vccd1 hold516/X sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_40_434 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_40_445 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_12_158 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
Xhold549 _0996_/X vssd1 vssd1 vccd1 vccd1 hold549/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold538 la_data_in[23] vssd1 vssd1 vccd1 vccd1 hold538/X sky130_fd_sc_hd__dlygate4sd3_1
XTAP_810 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_21_681 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_843 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_832 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_821 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_876 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_865 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_854 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_57_96 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_2315_ _2315_/CLK _2315_/D _2054_/Y vssd1 vssd1 vccd1 vccd1 _2315_/Q sky130_fd_sc_hd__dfrtp_1
XTAP_887 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_2246_ _2249_/CLK _2246_/D _1985_/Y vssd1 vssd1 vccd1 vccd1 _2246_/Q sky130_fd_sc_hd__dfrtp_1
XFILLER_0_18_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__1311__B1 _1541_/B1 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_2177_ _2177_/CLK _2177_/D _1917_/Y vssd1 vssd1 vccd1 vccd1 _2177_/Q sky130_fd_sc_hd__dfrtp_4
X_1128_ _2192_/Q _2100_/Q _1156_/S vssd1 vssd1 vccd1 vccd1 _1128_/X sky130_fd_sc_hd__mux2_1
XANTENNA__1679__A _2107_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_1059_ hold573/X _1097_/A2 _1097_/B1 _1058_/X vssd1 vssd1 vccd1 vccd1 _2315_/D sky130_fd_sc_hd__a22o_1
XFILLER_0_48_567 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__1614__A1 _2079_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_36_707 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_8_653 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xcontroller_624 vssd1 vssd1 vccd1 vccd1 controller_624/HI la_data_out[6] sky130_fd_sc_hd__conb_1
XFILLER_0_35_228 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA_fanout608_A _2034_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xcontroller_646 vssd1 vssd1 vccd1 vccd1 controller_646/HI la_data_out[28] sky130_fd_sc_hd__conb_1
Xcontroller_635 vssd1 vssd1 vccd1 vccd1 controller_635/HI la_data_out[17] sky130_fd_sc_hd__conb_1
Xcontroller_657 vssd1 vssd1 vccd1 vccd1 controller_657/HI la_data_out[121] sky130_fd_sc_hd__conb_1
XFILLER_0_31_401 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_31_445 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_3_391 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xinput136 data_in[75] vssd1 vssd1 vccd1 vccd1 _1481_/A1 sky130_fd_sc_hd__clkbuf_2
Xinput103 data_in[45] vssd1 vssd1 vccd1 vccd1 _1541_/A1 sky130_fd_sc_hd__buf_1
Xinput114 data_in[55] vssd1 vssd1 vccd1 vccd1 _1521_/A1 sky130_fd_sc_hd__buf_1
Xinput125 data_in[65] vssd1 vssd1 vccd1 vccd1 _1501_/A1 sky130_fd_sc_hd__clkbuf_2
Xinput158 data_in[95] vssd1 vssd1 vccd1 vccd1 _1407_/A1 sky130_fd_sc_hd__buf_1
Xinput147 data_in[85] vssd1 vssd1 vccd1 vccd1 _1437_/A1 sky130_fd_sc_hd__buf_1
Xinput169 hold83/X vssd1 vssd1 vccd1 vccd1 hold84/A sky130_fd_sc_hd__clkbuf_1
XANTENNA__1302__B1 _1527_/B1 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_39_512 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_39_534 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__1605__B2 _2084_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__1081__A2 _1095_/A2 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__1528__S hold80/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_41_209 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_34_294 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_128 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_139 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_2100_ _2182_/CLK _2100_/D _1843_/Y vssd1 vssd1 vccd1 vccd1 _2100_/Q sky130_fd_sc_hd__dfrtp_4
XANTENNA__1541__B1 _1541_/B1 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_2031_ _2033_/A vssd1 vssd1 vccd1 vccd1 _2031_/Y sky130_fd_sc_hd__inv_2
XFILLER_0_27_99 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XPHY_0 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_9_428 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_45_515 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_45_559 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_1815_ _1988_/A vssd1 vssd1 vccd1 vccd1 _1815_/Y sky130_fd_sc_hd__inv_2
XANTENNA__1438__S hold27/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_1746_ _2184_/Q _1756_/B vssd1 vssd1 vccd1 vccd1 _1746_/X sky130_fd_sc_hd__and2_1
Xhold302 hold902/X vssd1 vssd1 vccd1 vccd1 hold302/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold324 hold324/A vssd1 vssd1 vccd1 vccd1 _1250_/B sky130_fd_sc_hd__dlygate4sd3_1
Xhold335 hold335/A vssd1 vssd1 vccd1 vccd1 _1334_/B sky130_fd_sc_hd__dlygate4sd3_1
Xhold313 _1248_/X vssd1 vssd1 vccd1 vccd1 hold313/X sky130_fd_sc_hd__dlygate4sd3_1
X_1677_ _2105_/Q _1677_/B vssd1 vssd1 vccd1 vccd1 _1677_/X sky130_fd_sc_hd__and2_1
XANTENNA__1962__A _2002_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xhold368 hold368/A vssd1 vssd1 vccd1 vccd1 _1340_/B sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_7_76 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xhold346 hold362/X vssd1 vssd1 vccd1 vccd1 hold346/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold357 hold387/X vssd1 vssd1 vccd1 vccd1 hold357/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold379 _1244_/X vssd1 vssd1 vccd1 vccd1 hold379/X sky130_fd_sc_hd__buf_1
XTAP_651 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__1681__B _1725_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_640 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_695 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_684 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_673 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_662 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_fanout558_A _1023_/Y vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_2229_ _2322_/CLK _2229_/D _1969_/Y vssd1 vssd1 vccd1 vccd1 _2229_/Q sky130_fd_sc_hd__dfrtp_1
XANTENNA__1063__A2 _1097_/A2 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_36_559 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_44_592 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_16_283 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_31_253 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__1872__A _2002_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xhold880 _2275_/Q vssd1 vssd1 vccd1 vccd1 hold880/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold891 la_data_in[41] vssd1 vssd1 vccd1 vccd1 hold891/X sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA__1523__B1 _1527_/B1 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_hold937_A _2101_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_39_375 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_27_537 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_1600_ _1599_/X _2086_/Q _1622_/S vssd1 vssd1 vccd1 vccd1 _1600_/X sky130_fd_sc_hd__mux2_1
XANTENNA__1258__S hold26/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xoutput407 _1725_/X vssd1 vssd1 vccd1 vccd1 data_out[83] sky130_fd_sc_hd__buf_12
XFILLER_0_22_253 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
Xoutput418 _1735_/X vssd1 vssd1 vccd1 vccd1 data_out[93] sky130_fd_sc_hd__buf_12
XANTENNA__1782__A _2220_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_10_415 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xoutput429 hold594/X vssd1 vssd1 vccd1 vccd1 la_data_out[102] sky130_fd_sc_hd__buf_12
X_1531_ _1531_/A1 _1533_/A2 _1533_/B1 _2121_/Q hold164/X vssd1 vssd1 vccd1 vccd1 _1531_/X
+ sky130_fd_sc_hd__a221o_1
X_1462_ _1527_/A2 hold122/X _1022_/B _1277_/A vssd1 vssd1 vccd1 vccd1 _1462_/X sky130_fd_sc_hd__a211o_1
X_1393_ _1392_/X hold970/X _1435_/S vssd1 vssd1 vccd1 vccd1 _2180_/D sky130_fd_sc_hd__mux2_1
XFILLER_0_54_53 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_2014_ _2033_/A vssd1 vssd1 vccd1 vccd1 _2014_/Y sky130_fd_sc_hd__inv_2
XFILLER_0_9_214 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__1293__A2 _1529_/A2 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__1957__A _1957_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_18_504 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__1045__A2 _1095_/A2 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__1168__S _1188_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xhold110 _1002_/Y vssd1 vssd1 vccd1 vccd1 hold110/X sky130_fd_sc_hd__dlygate4sd3_1
X_1729_ _2167_/Q _1761_/B vssd1 vssd1 vccd1 vccd1 _1729_/X sky130_fd_sc_hd__and2_1
Xhold121 _1025_/Y vssd1 vssd1 vccd1 vccd1 _1198_/C sky130_fd_sc_hd__dlygate4sd3_1
Xhold132 _1400_/X vssd1 vssd1 vccd1 vccd1 hold132/X sky130_fd_sc_hd__dlymetal6s2s_1
Xhold143 _1303_/X vssd1 vssd1 vccd1 vccd1 _2210_/D sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA__1692__A _2120_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xhold154 hold216/X vssd1 vssd1 vccd1 vccd1 hold154/X sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_1_670 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
Xhold176 _1436_/X vssd1 vssd1 vccd1 vccd1 hold176/X sky130_fd_sc_hd__buf_1
Xhold165 _1296_/X vssd1 vssd1 vccd1 vccd1 hold165/X sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_1_681 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
Xfanout612 _2061_/A vssd1 vssd1 vccd1 vccd1 _2065_/A sky130_fd_sc_hd__buf_8
Xhold187 _1421_/X vssd1 vssd1 vccd1 vccd1 hold187/X sky130_fd_sc_hd__buf_1
Xhold198 _1314_/X vssd1 vssd1 vccd1 vccd1 hold198/X sky130_fd_sc_hd__dlygate4sd3_1
Xfanout601 _1922_/A vssd1 vssd1 vccd1 vccd1 _1916_/A sky130_fd_sc_hd__buf_8
XANTENNA__1505__B1 _1519_/B1 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_470 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_481 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_492 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__1284__A2 _1529_/A2 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_36_378 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_17_570 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_32_540 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_20_713 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__1275__A2 _1529_/A2 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_24_45 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__1777__A _2215_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_0962_ _0992_/A _0992_/B vssd1 vssd1 vccd1 vccd1 _0978_/B sky130_fd_sc_hd__or2_2
XFILLER_0_40_66 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_2_401 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_40_99 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_1514_ hold464/X _2129_/Q _1520_/S vssd1 vssd1 vccd1 vccd1 _1514_/X sky130_fd_sc_hd__mux2_1
XFILLER_0_49_75 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_1445_ _1445_/A hold48/X vssd1 vssd1 vccd1 vccd1 hold49/A sky130_fd_sc_hd__and2_1
X_1376_ _1394_/A _1376_/B vssd1 vssd1 vccd1 vccd1 _1376_/X sky130_fd_sc_hd__and2_1
XANTENNA__1266__A2 _1519_/A2 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_37_109 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__1687__A _2115_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_18_378 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_18_389 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__1257__A2 _1519_/A2 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_37_676 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_24_304 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_36_186 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_36_197 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_51_189 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_51_167 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__1536__S hold80/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_1230_ input61/X _1503_/A2 _1503_/B1 _2235_/Q hold348/X vssd1 vssd1 vccd1 vccd1 _1230_/X
+ sky130_fd_sc_hd__a221o_1
X_1161_ _2264_/Q _1189_/A2 _1189_/B1 _1160_/X vssd1 vssd1 vccd1 vccd1 _1161_/X sky130_fd_sc_hd__a22o_1
Xclkbuf_leaf_26_wb_clk_i clkbuf_leaf_9_wb_clk_i/A vssd1 vssd1 vccd1 vccd1 _2164_/CLK
+ sky130_fd_sc_hd__clkbuf_16
X_1092_ _2210_/Q _2118_/Q _1188_/S vssd1 vssd1 vccd1 vccd1 _1092_/X sky130_fd_sc_hd__mux2_1
XFILLER_0_35_66 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_51_54 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_1994_ _2008_/A vssd1 vssd1 vccd1 vccd1 _1994_/Y sky130_fd_sc_hd__inv_2
XFILLER_0_42_101 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_15_326 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_42_145 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_42_123 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_15_337 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_2_253 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_2_264 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__1184__A1 _2072_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__1970__A _1979_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_48_3 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_1428_ _1428_/A1 _1569_/A2 _1569_/B1 _2169_/Q hold64/X vssd1 vssd1 vccd1 vccd1 hold65/A
+ sky130_fd_sc_hd__a221o_1
X_1359_ input14/X _1529_/A2 _1529_/B1 _2192_/Q hold290/X vssd1 vssd1 vccd1 vccd1 _1359_/X
+ sky130_fd_sc_hd__a221o_1
XANTENNA__1487__A2 _1503_/A2 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout540_A _1724_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_38_429 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_46_462 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_18_164 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__1880__A _2069_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_24_101 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_37_473 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XANTENNA_output292_A _1768_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_21_57 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_12_307 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xhold709 hold905/X vssd1 vssd1 vccd1 vccd1 hold709/X sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_24_167 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_40_638 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__1166__A1 _2081_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_20_362 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_2262_ _2296_/CLK _2262_/D _2001_/Y vssd1 vssd1 vccd1 vccd1 _2262_/Q sky130_fd_sc_hd__dfrtp_1
X_1213_ _1212_/X _2240_/Q _1252_/S vssd1 vssd1 vccd1 vccd1 _1213_/X sky130_fd_sc_hd__mux2_1
X_2193_ _2217_/CLK _2193_/D _1933_/Y vssd1 vssd1 vccd1 vccd1 _2193_/Q sky130_fd_sc_hd__dfrtp_4
XANTENNA__1469__A2 _1197_/D vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_1144_ _2184_/Q _2092_/Q _1156_/S vssd1 vssd1 vccd1 vccd1 _1144_/X sky130_fd_sc_hd__mux2_1
X_1075_ hold636/X _1095_/A2 _1095_/B1 _1074_/X vssd1 vssd1 vccd1 vccd1 _2307_/D sky130_fd_sc_hd__a22o_1
XFILLER_0_7_312 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_16_635 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_28_473 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_1977_ _1979_/A vssd1 vssd1 vccd1 vccd1 _1977_/Y sky130_fd_sc_hd__inv_2
XFILLER_0_16_657 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__1965__A _2026_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_43_465 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__1684__B _1725_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_24_690 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_30_148 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA_fanout588_A _1038_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xhold14 hold14/A vssd1 vssd1 vccd1 vccd1 hold14/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold36 hold36/A vssd1 vssd1 vccd1 vccd1 hold36/X sky130_fd_sc_hd__dlymetal6s2s_1
Xhold47 hold47/A vssd1 vssd1 vccd1 vccd1 hold47/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold25 hold39/X vssd1 vssd1 vccd1 vccd1 hold40/A sky130_fd_sc_hd__dlygate4sd3_1
Xhold69 hold69/A vssd1 vssd1 vccd1 vccd1 hold69/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold58 hold58/A vssd1 vssd1 vccd1 vccd1 hold58/X sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA__1617__C1 hold117/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__2036__A _2065_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__1093__B1 _1097_/B1 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_38_259 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__1875__A _2002_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_34_454 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_34_465 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_21_137 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__1148__A1 _2090_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_hold967_A _2167_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_30_660 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_16_13 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_16_57 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__1320__A1 input28/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__1320__B2 _2205_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_29_237 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_1900_ _1913_/A vssd1 vssd1 vccd1 vccd1 _1900_/Y sky130_fd_sc_hd__inv_2
XANTENNA__1623__A2 _1623_/A2 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__1084__A0 _2214_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_1831_ _1852_/A vssd1 vssd1 vccd1 vccd1 _1831_/Y sky130_fd_sc_hd__inv_2
XFILLER_0_44_218 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__1785__A _2223_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_37_281 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_1762_ _2200_/Q _1766_/B vssd1 vssd1 vccd1 vccd1 _1762_/X sky130_fd_sc_hd__and2_1
Xhold506 _1512_/X vssd1 vssd1 vccd1 vccd1 _2130_/D sky130_fd_sc_hd__dlygate4sd3_1
Xhold517 la_data_in[75] vssd1 vssd1 vccd1 vccd1 hold517/X sky130_fd_sc_hd__dlygate4sd3_1
X_1693_ _2121_/Q _1715_/B vssd1 vssd1 vccd1 vccd1 _1693_/X sky130_fd_sc_hd__and2_1
Xhold528 _1808_/D vssd1 vssd1 vccd1 vccd1 _1382_/B sky130_fd_sc_hd__dlygate4sd3_1
Xhold539 la_data_in[86] vssd1 vssd1 vccd1 vccd1 hold539/X sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_40_457 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_800 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_21_671 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_57_53 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_844 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_833 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_822 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_811 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_877 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_866 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_855 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_2314_ _2330_/CLK _2314_/D _2053_/Y vssd1 vssd1 vccd1 vccd1 _2314_/Q sky130_fd_sc_hd__dfrtp_1
XTAP_888 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_2245_ _2249_/CLK _2245_/D _1984_/Y vssd1 vssd1 vccd1 vccd1 _2245_/Q sky130_fd_sc_hd__dfrtp_1
X_2176_ _2177_/CLK _2176_/D _1916_/Y vssd1 vssd1 vccd1 vccd1 _2176_/Q sky130_fd_sc_hd__dfrtp_4
X_1127_ hold615/X _1189_/A2 _1189_/B1 _1126_/X vssd1 vssd1 vccd1 vccd1 _2281_/D sky130_fd_sc_hd__a22o_1
XANTENNA__1311__B2 _2208_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_clkbuf_leaf_2_wb_clk_i_A clkbuf_leaf_9_wb_clk_i/A vssd1 vssd1 vccd1 vccd1
+ sky130_fd_sc_hd__diode_2
XFILLER_0_48_513 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_1058_ _2227_/Q _2135_/Q _1094_/S vssd1 vssd1 vccd1 vccd1 _1058_/X sky130_fd_sc_hd__mux2_1
XFILLER_0_8_621 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__1075__B1 _1095_/B1 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_8_643 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__1695__A _2123_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xcontroller_625 vssd1 vssd1 vccd1 vccd1 controller_625/HI la_data_out[7] sky130_fd_sc_hd__conb_1
Xcontroller_636 vssd1 vssd1 vccd1 vccd1 controller_636/HI la_data_out[18] sky130_fd_sc_hd__conb_1
Xcontroller_647 vssd1 vssd1 vccd1 vccd1 controller_647/HI la_data_out[29] sky130_fd_sc_hd__conb_1
XFILLER_0_16_432 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_43_284 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xinput115 data_in[56] vssd1 vssd1 vccd1 vccd1 _1519_/A1 sky130_fd_sc_hd__buf_1
Xinput104 data_in[46] vssd1 vssd1 vccd1 vccd1 _1539_/A1 sky130_fd_sc_hd__dlymetal6s2s_1
Xinput126 data_in[66] vssd1 vssd1 vccd1 vccd1 _1499_/A1 sky130_fd_sc_hd__clkbuf_2
Xinput159 data_in[96] vssd1 vssd1 vccd1 vccd1 _1404_/A1 sky130_fd_sc_hd__buf_1
Xinput148 data_in[86] vssd1 vssd1 vccd1 vccd1 _1434_/A1 sky130_fd_sc_hd__buf_1
Xinput137 data_in[76] vssd1 vssd1 vccd1 vccd1 _1479_/A1 sky130_fd_sc_hd__clkbuf_2
XANTENNA__1302__B2 _2211_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XPHY_110 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__1066__A0 _2223_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__1605__A2 _1623_/A2 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__1369__A1 _2188_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_22_402 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_129 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__1544__S hold80/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__1541__A1 _1541_/A1 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__1541__B2 _2116_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_27_23 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_2030_ _2033_/A vssd1 vssd1 vccd1 vccd1 _2030_/Y sky130_fd_sc_hd__inv_2
XFILLER_0_9_407 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XPHY_1 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_43_99 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_43_77 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_45_505 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_1814_ _1988_/A vssd1 vssd1 vccd1 vccd1 _1814_/Y sky130_fd_sc_hd__inv_2
XFILLER_0_25_240 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_1745_ _2183_/Q _1756_/B vssd1 vssd1 vccd1 vccd1 _1745_/X sky130_fd_sc_hd__and2_1
Xhold303 la_data_in[77] vssd1 vssd1 vccd1 vccd1 hold303/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold325 _1250_/X vssd1 vssd1 vccd1 vccd1 hold325/X sky130_fd_sc_hd__buf_1
Xhold314 _1249_/X vssd1 vssd1 vccd1 vccd1 _2228_/D sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_40_232 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_1676_ _2104_/Q _1677_/B vssd1 vssd1 vccd1 vccd1 _1676_/X sky130_fd_sc_hd__and2_1
Xhold358 hold358/A vssd1 vssd1 vccd1 vccd1 _1241_/B sky130_fd_sc_hd__dlygate4sd3_1
Xhold347 hold347/A vssd1 vssd1 vccd1 vccd1 _1229_/B sky130_fd_sc_hd__dlygate4sd3_1
Xhold336 _1334_/X vssd1 vssd1 vccd1 vccd1 hold336/X sky130_fd_sc_hd__buf_1
Xhold369 _1340_/X vssd1 vssd1 vccd1 vccd1 hold369/X sky130_fd_sc_hd__buf_1
XTAP_652 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_641 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_630 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_685 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_674 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_663 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__1532__A1 _2120_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_696 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_30_3 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_2228_ _2322_/CLK _2228_/D _1968_/Y vssd1 vssd1 vccd1 vccd1 _2228_/Q sky130_fd_sc_hd__dfrtp_1
X_2159_ _2249_/CLK hold91/X _1900_/Y vssd1 vssd1 vccd1 vccd1 _2159_/Q sky130_fd_sc_hd__dfrtp_1
XANTENNA__1296__B1 _1529_/B1 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_48_343 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XANTENNA__1599__B2 _2087_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_36_516 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_8_473 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_44_582 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_31_210 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
Xhold881 la_data_in[42] vssd1 vssd1 vccd1 vccd1 hold881/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold870 _1327_/X vssd1 vssd1 vccd1 vccd1 _2202_/D sky130_fd_sc_hd__dlygate4sd3_1
Xhold892 _1324_/X vssd1 vssd1 vccd1 vccd1 _2203_/D sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA__1523__B2 _2125_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__1287__B1 _1529_/B1 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_39_332 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_54_302 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_54_379 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_23_700 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
Xoutput408 _1726_/X vssd1 vssd1 vccd1 vccd1 data_out[84] sky130_fd_sc_hd__buf_12
Xoutput419 _1736_/X vssd1 vssd1 vccd1 vccd1 data_out[94] sky130_fd_sc_hd__buf_12
XFILLER_0_22_265 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_1530_ _1529_/X _2121_/Q _1530_/S vssd1 vssd1 vccd1 vccd1 _1530_/X sky130_fd_sc_hd__mux2_1
X_1461_ hold123/X _2157_/Q _1461_/S vssd1 vssd1 vccd1 vccd1 _1461_/X sky130_fd_sc_hd__mux2_1
X_1392_ input2/X _1569_/A2 _1569_/B1 _2181_/Q _1391_/X vssd1 vssd1 vccd1 vccd1 _1392_/X
+ sky130_fd_sc_hd__a221o_1
XFILLER_0_38_33 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_54_21 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__1278__B1 _1519_/B1 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_2013_ _2033_/A vssd1 vssd1 vccd1 vccd1 _2013_/Y sky130_fd_sc_hd__inv_2
XFILLER_0_54_76 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_45_335 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__1450__B1 _1545_/B1 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__1973__A _1979_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xhold100 hold100/A vssd1 vssd1 vccd1 vccd1 _1418_/B sky130_fd_sc_hd__dlygate4sd3_1
Xhold133 _1401_/X vssd1 vssd1 vccd1 vccd1 hold133/X sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_41_585 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xhold122 _1027_/Y vssd1 vssd1 vccd1 vccd1 hold122/X sky130_fd_sc_hd__clkdlybuf4s25_1
Xhold111 _1459_/Y vssd1 vssd1 vccd1 vccd1 hold111/X sky130_fd_sc_hd__clkdlybuf4s25_1
Xhold144 la_data_in[33] vssd1 vssd1 vccd1 vccd1 hold144/X sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA__1202__B1 _1193_/Y vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_13_276 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_1728_ _2166_/Q _1761_/B vssd1 vssd1 vccd1 vccd1 _1728_/X sky130_fd_sc_hd__and2_1
X_1659_ _2087_/Q _1677_/B vssd1 vssd1 vccd1 vccd1 _1659_/X sky130_fd_sc_hd__and2_1
Xhold155 hold155/A vssd1 vssd1 vccd1 vccd1 _1412_/B sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA__1184__S _1188_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xhold177 _1625_/X vssd1 vssd1 vccd1 vccd1 hold177/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold166 _1297_/X vssd1 vssd1 vccd1 vccd1 _2212_/D sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA__1692__B _1715_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xhold199 la_data_in[46] vssd1 vssd1 vccd1 vccd1 hold57/A sky130_fd_sc_hd__dlygate4sd3_1
Xfanout613 _2061_/A vssd1 vssd1 vccd1 vccd1 _2069_/A sky130_fd_sc_hd__buf_8
Xhold188 _1615_/X vssd1 vssd1 vccd1 vccd1 hold188/X sky130_fd_sc_hd__dlygate4sd3_1
Xfanout602 input262/X vssd1 vssd1 vccd1 vccd1 _1922_/A sky130_fd_sc_hd__buf_8
XANTENNA__1505__A1 _1505_/A1 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_460 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_fanout570_A _1519_/A2 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_471 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_482 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_493 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__1269__B1 _1519_/B1 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_48_173 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_8_281 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__2044__A _2065_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__1883__A _1979_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__1094__S _1094_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_32_596 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_59_449 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_24_79 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_39_151 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_55_633 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_0961_ hold76/X _1014_/B hold21/X _1002_/A vssd1 vssd1 vccd1 vccd1 _0978_/A sky130_fd_sc_hd__or4_2
XFILLER_0_42_305 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_40_78 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_23_530 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_23_541 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_35_390 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_50_360 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_1513_ _1513_/A1 _1519_/A2 _1519_/B1 _2130_/Q hold463/X vssd1 vssd1 vccd1 vccd1 _1513_/X
+ sky130_fd_sc_hd__a221o_1
XFILLER_0_23_596 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_1444_ _1443_/X _2163_/Q hold27/X vssd1 vssd1 vccd1 vccd1 hold41/A sky130_fd_sc_hd__mux2_1
X_1375_ hold128/X _2186_/Q _1435_/S vssd1 vssd1 vccd1 vccd1 _1375_/X sky130_fd_sc_hd__mux2_1
XFILLER_0_4_78 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__1687__B _1724_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_18_346 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_18_368 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_41_393 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_290 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__2039__A _2039_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__1878__A _2039_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_49_460 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_37_655 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_51_113 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_51_124 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_20_533 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_19_57 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_1160_ _2176_/Q _2084_/Q _1178_/S vssd1 vssd1 vccd1 vccd1 _1160_/X sky130_fd_sc_hd__mux2_1
XANTENNA__1350__C1 hold406/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_1091_ hold574/X _1097_/A2 _1097_/B1 _1090_/X vssd1 vssd1 vccd1 vccd1 _2299_/D sky130_fd_sc_hd__a22o_1
XFILLER_0_35_45 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_59_279 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_7_505 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_1993_ _2008_/A vssd1 vssd1 vccd1 vccd1 _1993_/Y sky130_fd_sc_hd__inv_2
XFILLER_0_43_625 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_27_154 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_27_165 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_1427_ _1445_/A hold63/X vssd1 vssd1 vccd1 vccd1 hold64/A sky130_fd_sc_hd__and2_1
X_1358_ _1415_/A _1358_/B vssd1 vssd1 vccd1 vccd1 _1358_/X sky130_fd_sc_hd__and2_1
X_1289_ _1310_/A _1289_/B vssd1 vssd1 vccd1 vccd1 _1289_/X sky130_fd_sc_hd__and2_1
XANTENNA__1698__A _2126_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_19_655 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_19_666 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_34_636 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_33_113 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__1175__A2 _1189_/A2 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_37_430 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_21_36 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_25_603 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_25_625 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_37_485 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_20_341 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_2330_ _2330_/CLK _2330_/D _2069_/Y vssd1 vssd1 vccd1 vccd1 _2330_/Q sky130_fd_sc_hd__dfrtp_1
XANTENNA__1571__C1 hold276/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_2261_ _2269_/CLK _2261_/D _2000_/Y vssd1 vssd1 vccd1 vccd1 _2261_/Q sky130_fd_sc_hd__dfrtp_1
XANTENNA__1282__S hold26/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_1212_ input68/X _1463_/B _1499_/B1 _2241_/Q hold231/X vssd1 vssd1 vccd1 vccd1 _1212_/X
+ sky130_fd_sc_hd__a221o_1
X_2192_ _2194_/CLK _2192_/D _1932_/Y vssd1 vssd1 vccd1 vccd1 _2192_/Q sky130_fd_sc_hd__dfrtp_4
X_1143_ hold616/X _1189_/A2 _1189_/B1 _1142_/X vssd1 vssd1 vccd1 vccd1 _2273_/D sky130_fd_sc_hd__a22o_1
X_1074_ _2219_/Q _2127_/Q _1086_/S vssd1 vssd1 vccd1 vccd1 _1074_/X sky130_fd_sc_hd__mux2_1
XFILLER_0_47_205 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_1_79 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_1_68 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_47_216 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_47_249 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_1976_ _1979_/A vssd1 vssd1 vccd1 vccd1 _1976_/Y sky130_fd_sc_hd__inv_2
XFILLER_0_43_422 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_15_113 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_43_477 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_31_617 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XANTENNA__1157__A2 _1157_/A2 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xhold15 hold15/A vssd1 vssd1 vccd1 vccd1 hold15/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold37 hold37/A vssd1 vssd1 vccd1 vccd1 hold37/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold26 hold26/A vssd1 vssd1 vccd1 vccd1 hold26/X sky130_fd_sc_hd__buf_8
Xhold48 hold48/A vssd1 vssd1 vccd1 vccd1 hold48/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold59 hold59/A vssd1 vssd1 vccd1 vccd1 hold59/X sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_19_463 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_34_477 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_21_127 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_30_672 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__1320__A2 _1527_/A2 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_57_558 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_1830_ _1852_/A vssd1 vssd1 vccd1 vccd1 _1830_/Y sky130_fd_sc_hd__inv_2
X_1761_ _2199_/Q _1761_/B vssd1 vssd1 vccd1 vccd1 _1761_/X sky130_fd_sc_hd__and2_1
XFILLER_0_4_327 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
Xhold518 _1222_/X vssd1 vssd1 vccd1 vccd1 _2237_/D sky130_fd_sc_hd__dlygate4sd3_1
Xhold507 la_data_in[17] vssd1 vssd1 vccd1 vccd1 hold507/X sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_25_499 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_1692_ _2120_/Q _1715_/B vssd1 vssd1 vccd1 vccd1 _1692_/X sky130_fd_sc_hd__and2_1
Xhold529 _1382_/X vssd1 vssd1 vccd1 vccd1 hold529/X sky130_fd_sc_hd__dlymetal6s2s_1
XTAP_801 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_20_160 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_834 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_823 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_812 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_2313_ _2315_/CLK _2313_/D _2052_/Y vssd1 vssd1 vccd1 vccd1 _2313_/Q sky130_fd_sc_hd__dfrtp_1
XTAP_867 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_856 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_845 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_889 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_878 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_2244_ _2249_/CLK hold4/X _1983_/Y vssd1 vssd1 vccd1 vccd1 _2244_/Q sky130_fd_sc_hd__dfrtp_1
Xclkbuf_leaf_10_wb_clk_i clkbuf_1_1__f_wb_clk_i/X vssd1 vssd1 vccd1 vccd1 _2225_/CLK
+ sky130_fd_sc_hd__clkbuf_16
X_2175_ _2177_/CLK _2175_/D _1915_/Y vssd1 vssd1 vccd1 vccd1 _2175_/Q sky130_fd_sc_hd__dfrtp_4
X_1126_ _2193_/Q _2101_/Q _1156_/S vssd1 vssd1 vccd1 vccd1 _1126_/X sky130_fd_sc_hd__mux2_1
XANTENNA__1311__A2 _1197_/D vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_1057_ hold589/X _1057_/A2 _1057_/B1 _1056_/X vssd1 vssd1 vccd1 vccd1 _2316_/D sky130_fd_sc_hd__a22o_1
XANTENNA__1075__B2 _1074_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_16_400 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__1976__A _1979_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__1695__B _1715_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xcontroller_626 vssd1 vssd1 vccd1 vccd1 controller_626/HI la_data_out[8] sky130_fd_sc_hd__conb_1
Xcontroller_637 vssd1 vssd1 vccd1 vccd1 controller_637/HI la_data_out[19] sky130_fd_sc_hd__conb_1
Xcontroller_648 vssd1 vssd1 vccd1 vccd1 controller_648/HI la_data_out[30] sky130_fd_sc_hd__conb_1
XFILLER_0_16_444 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_16_477 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_1959_ _2002_/A vssd1 vssd1 vccd1 vccd1 _1959_/Y sky130_fd_sc_hd__inv_2
XFILLER_0_3_393 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_12_661 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xinput116 data_in[57] vssd1 vssd1 vccd1 vccd1 _1517_/A1 sky130_fd_sc_hd__buf_1
Xinput105 data_in[47] vssd1 vssd1 vccd1 vccd1 _1537_/A1 sky130_fd_sc_hd__buf_1
Xinput127 data_in[67] vssd1 vssd1 vccd1 vccd1 _1497_/A1 sky130_fd_sc_hd__buf_2
Xinput138 data_in[77] vssd1 vssd1 vccd1 vccd1 _1477_/A1 sky130_fd_sc_hd__buf_2
Xinput149 data_in[87] vssd1 vssd1 vccd1 vccd1 _1431_/A1 sky130_fd_sc_hd__buf_1
XANTENNA_hold276_A _1355_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__1302__A2 _1197_/D vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_hold443_A _1223_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XPHY_100 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__2047__A _2065_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_39_503 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XPHY_111 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_26_208 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__1886__A _1979_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_22_414 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_22_447 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__1541__A2 _1197_/D vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_27_57 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_27_68 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_43_45 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XPHY_2 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_45_528 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_38_580 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_1813_ _2249_/Q vssd1 vssd1 vccd1 vccd1 _1813_/X sky130_fd_sc_hd__clkbuf_1
X_1744_ _2182_/Q _1756_/B vssd1 vssd1 vccd1 vccd1 _1744_/X sky130_fd_sc_hd__and2_1
XFILLER_0_40_200 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xhold304 _1216_/X vssd1 vssd1 vccd1 vccd1 _2239_/D sky130_fd_sc_hd__dlygate4sd3_1
Xhold315 hold321/X vssd1 vssd1 vccd1 vccd1 hold315/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold326 _1251_/X vssd1 vssd1 vccd1 vccd1 hold326/X sky130_fd_sc_hd__dlygate4sd3_1
X_1675_ _2103_/Q _1677_/B vssd1 vssd1 vccd1 vccd1 _1675_/X sky130_fd_sc_hd__and2_1
Xhold359 _1241_/X vssd1 vssd1 vccd1 vccd1 hold359/X sky130_fd_sc_hd__buf_1
Xhold348 _1229_/X vssd1 vssd1 vccd1 vccd1 hold348/X sky130_fd_sc_hd__clkbuf_2
Xhold337 _1335_/X vssd1 vssd1 vccd1 vccd1 hold337/X sky130_fd_sc_hd__dlygate4sd3_1
XTAP_620 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_642 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_631 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_686 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_675 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_664 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_653 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_697 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_2227_ _2239_/CLK _2227_/D _1967_/Y vssd1 vssd1 vccd1 vccd1 _2227_/Q sky130_fd_sc_hd__dfrtp_1
XANTENNA__1470__S hold80/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_23_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_2158_ _2251_/CLK _2158_/D _1899_/Y vssd1 vssd1 vccd1 vccd1 _2158_/Q sky130_fd_sc_hd__dfrtp_1
XANTENNA__1296__B2 _2213_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_2089_ _2182_/CLK _2089_/D _1832_/Y vssd1 vssd1 vccd1 vccd1 _2089_/Q sky130_fd_sc_hd__dfrtp_4
XFILLER_0_48_300 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_1109_ _2290_/Q _1139_/A2 _1139_/B1 _1108_/X vssd1 vssd1 vccd1 vccd1 _1109_/X sky130_fd_sc_hd__a22o_1
XFILLER_0_48_388 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_48_355 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_16_241 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_32_712 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
Xhold860 _2152_/Q vssd1 vssd1 vccd1 vccd1 hold860/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold871 _2301_/Q vssd1 vssd1 vccd1 vccd1 hold871/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold882 _1548_/X vssd1 vssd1 vccd1 vccd1 _2112_/D sky130_fd_sc_hd__dlygate4sd3_1
Xhold893 _2294_/Q vssd1 vssd1 vccd1 vccd1 hold893/X sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA__1523__A2 _1527_/A2 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__1287__B2 _2216_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__1039__B2 _1038_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_39_399 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_23_712 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_35_572 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_50_520 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xoutput409 _1727_/X vssd1 vssd1 vccd1 vccd1 data_out[85] sky130_fd_sc_hd__buf_12
XANTENNA_output365_A _1687_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_1460_ _1527_/A2 hold122/X _1541_/B1 hold111/X vssd1 vssd1 vccd1 vccd1 _1460_/X sky130_fd_sc_hd__a211o_1
XFILLER_0_22_299 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_1391_ _1394_/A hold88/X vssd1 vssd1 vccd1 vccd1 _1391_/X sky130_fd_sc_hd__and2_2
XFILLER_0_38_45 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XANTENNA__1278__B2 _2219_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_2012_ _2033_/A vssd1 vssd1 vccd1 vccd1 _2012_/Y sky130_fd_sc_hd__inv_2
XFILLER_0_58_642 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_14_701 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
Xhold101 _1418_/X vssd1 vssd1 vccd1 vccd1 hold101/X sky130_fd_sc_hd__buf_1
XFILLER_0_41_575 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xhold123 _1460_/X vssd1 vssd1 vccd1 vccd1 hold123/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold134 hold153/X vssd1 vssd1 vccd1 vccd1 hold134/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold112 _1467_/X vssd1 vssd1 vccd1 vccd1 hold79/A sky130_fd_sc_hd__dlygate4sd3_1
X_1727_ _2165_/Q _1766_/B vssd1 vssd1 vccd1 vccd1 _1727_/X sky130_fd_sc_hd__and2_1
X_1658_ _2086_/Q _1680_/B vssd1 vssd1 vccd1 vccd1 _1658_/X sky130_fd_sc_hd__and2_1
XFILLER_0_41_597 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
Xhold145 hold257/X vssd1 vssd1 vccd1 vccd1 hold145/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold167 hold214/X vssd1 vssd1 vccd1 vccd1 hold167/X sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_13_288 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
Xhold156 _1412_/X vssd1 vssd1 vccd1 vccd1 hold156/X sky130_fd_sc_hd__buf_1
Xhold178 la_data_in[50] vssd1 vssd1 vccd1 vccd1 hold178/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold189 hold194/X vssd1 vssd1 vccd1 vccd1 hold189/X sky130_fd_sc_hd__dlygate4sd3_1
Xfanout614 _2061_/A vssd1 vssd1 vccd1 vccd1 _1982_/A sky130_fd_sc_hd__buf_4
Xfanout603 _1957_/A vssd1 vssd1 vccd1 vccd1 _1941_/A sky130_fd_sc_hd__buf_8
X_1589_ input77/X _1623_/A2 _1619_/B1 _2092_/Q hold529/X vssd1 vssd1 vccd1 vccd1 _1589_/X
+ sky130_fd_sc_hd__a221o_1
XANTENNA__1505__A2 _1519_/A2 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_450 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_472 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_461 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_483 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_494 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_fanout563_A _1003_/Y vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__1269__B2 _2222_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_48_141 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__1441__A1 _2164_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_24_509 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__1375__S _1435_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_hold775_A _2178_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__2060__A _2069_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xhold690 hold825/X vssd1 vssd1 vccd1 vccd1 hold690/X sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA_hold942_A _2085_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_clkbuf_leaf_26_wb_clk_i_A clkbuf_leaf_9_wb_clk_i/A vssd1 vssd1 vccd1 vccd1
+ sky130_fd_sc_hd__diode_2
X_0960_ hold76/X _1014_/B hold21/X _1002_/A vssd1 vssd1 vccd1 vccd1 _0990_/A sky130_fd_sc_hd__nor4_1
XFILLER_0_27_303 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_39_163 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_55_678 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_54_155 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_54_144 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_54_133 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_54_177 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_54_166 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_35_380 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__1285__S _1318_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_1512_ _1511_/X _2130_/Q _1520_/S vssd1 vssd1 vccd1 vccd1 _1512_/X sky130_fd_sc_hd__mux2_1
XFILLER_0_49_55 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_1443_ _1443_/A1 _1198_/A _1545_/B1 _2164_/Q hold31/X vssd1 vssd1 vccd1 vccd1 _1443_/X
+ sky130_fd_sc_hd__a221o_1
XANTENNA__1499__A1 _1499_/A1 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_1374_ input8/X _1533_/A2 _1533_/B1 _2187_/Q hold127/X vssd1 vssd1 vccd1 vccd1 _1374_/X
+ sky130_fd_sc_hd__a221o_1
XANTENNA__1120__A0 _2196_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_18_314 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_46_645 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__1423__A1 _2170_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_45_166 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_33_317 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_5_241 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_14_542 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__1187__B1 _1189_/B1 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_280 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_291 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_49_472 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__2055__A _2069_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_37_623 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__1414__A1 _2173_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__1894__A _1949_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_51_136 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_51_169 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XANTENNA__1178__A0 _2167_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_20_512 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_32_361 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_20_589 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_1090_ hold787/X _2119_/Q _1094_/S vssd1 vssd1 vccd1 vccd1 _1090_/X sky130_fd_sc_hd__mux2_1
XFILLER_0_35_57 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__1102__A0 _2205_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_51_34 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_1992_ _2008_/A vssd1 vssd1 vccd1 vccd1 _1992_/Y sky130_fd_sc_hd__inv_2
XFILLER_0_43_615 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_43_604 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_43_648 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_43_637 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_27_188 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_27_199 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_30_309 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_51_670 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_11_501 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__1169__B1 _1183_/B1 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_1426_ hold118/X hold977/X _1435_/S vssd1 vssd1 vccd1 vccd1 _2169_/D sky130_fd_sc_hd__mux2_1
X_1357_ hold277/X hold944/X _1372_/S vssd1 vssd1 vccd1 vccd1 _2192_/D sky130_fd_sc_hd__mux2_1
X_1288_ hold354/X _2215_/Q _1318_/S vssd1 vssd1 vccd1 vccd1 _1288_/X sky130_fd_sc_hd__mux2_1
XANTENNA__1979__A _1979_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__1698__B _1715_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_46_442 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_21_309 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_33_169 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_41_191 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__1332__B1 _1541_/B1 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__1889__A _2039_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__1194__C_N _1193_/Y vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_37_442 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_52_401 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_21_15 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_25_615 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_21_48 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_37_497 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_12_309 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_33_681 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__1571__B1 _1623_/B1 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_2260_ _2269_/CLK _2260_/D _1999_/Y vssd1 vssd1 vccd1 vccd1 _2260_/Q sky130_fd_sc_hd__dfrtp_1
X_1211_ _1277_/A _1211_/B vssd1 vssd1 vccd1 vccd1 _1211_/X sky130_fd_sc_hd__and2_1
X_2191_ _2194_/CLK _2191_/D _1931_/Y vssd1 vssd1 vccd1 vccd1 _2191_/Q sky130_fd_sc_hd__dfrtp_4
XANTENNA__1323__B1 _1541_/B1 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_1142_ _2185_/Q _2093_/Q _1178_/S vssd1 vssd1 vccd1 vccd1 _1142_/X sky130_fd_sc_hd__mux2_1
X_1073_ hold645/X _1095_/A2 _1095_/B1 _1072_/X vssd1 vssd1 vccd1 vccd1 _2308_/D sky130_fd_sc_hd__a22o_1
XFILLER_0_47_228 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_1975_ _1979_/A vssd1 vssd1 vccd1 vccd1 _1975_/Y sky130_fd_sc_hd__inv_2
XFILLER_0_16_626 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_28_464 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_43_434 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_15_136 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_16_648 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_28_497 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_15_158 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_31_629 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_53_3 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
Xhold16 hold16/A vssd1 vssd1 vccd1 vccd1 hold16/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold38 hold38/A vssd1 vssd1 vccd1 vccd1 hold38/X sky130_fd_sc_hd__clkbuf_2
X_1409_ _1415_/A _1409_/B vssd1 vssd1 vccd1 vccd1 _1409_/X sky130_fd_sc_hd__and2_1
Xhold27 hold27/A vssd1 vssd1 vccd1 vccd1 hold27/X sky130_fd_sc_hd__clkbuf_8
Xhold49 hold49/A vssd1 vssd1 vccd1 vccd1 hold49/X sky130_fd_sc_hd__buf_1
XANTENNA__1314__B1 _1527_/B1 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__1617__B2 _2078_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_38_217 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_38_228 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__1093__A2 _1097_/A2 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_53_209 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_46_272 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_19_486 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_22_607 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_15_681 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_21_106 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__1305__B1 _1541_/B1 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__1412__A _1415_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_29_206 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_25_401 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_1760_ _2198_/Q _1761_/B vssd1 vssd1 vccd1 vccd1 _1760_/X sky130_fd_sc_hd__and2_1
XFILLER_0_25_412 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_52_253 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_52_242 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
Xhold508 hold508/A vssd1 vssd1 vccd1 vccd1 hold508/X sky130_fd_sc_hd__dlygate4sd3_1
X_1691_ _2119_/Q _1724_/B vssd1 vssd1 vccd1 vccd1 _1691_/X sky130_fd_sc_hd__and2_1
Xhold519 hold531/X vssd1 vssd1 vccd1 vccd1 hold519/X sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_21_662 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_21_673 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_57_11 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_835 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_824 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_813 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_802 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_2312_ _2312_/CLK _2312_/D _2051_/Y vssd1 vssd1 vccd1 vccd1 _2312_/Q sky130_fd_sc_hd__dfrtp_1
XTAP_868 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_857 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_846 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_879 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_57_99 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_2243_ _2243_/D _1635_/C vssd1 vssd1 vccd1 vccd1 _2243_/Q sky130_fd_sc_hd__dlxtn_1
X_2174_ _2177_/CLK _2174_/D _1914_/Y vssd1 vssd1 vccd1 vccd1 _2174_/Q sky130_fd_sc_hd__dfrtp_4
X_1125_ hold642/X _1183_/A2 _1183_/B1 _1124_/X vssd1 vssd1 vccd1 vccd1 _2282_/D sky130_fd_sc_hd__a22o_1
X_1056_ _2228_/Q _2136_/Q _1094_/S vssd1 vssd1 vccd1 vccd1 _1056_/X sky130_fd_sc_hd__mux2_1
XANTENNA__1075__A2 _1095_/A2 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xcontroller_627 vssd1 vssd1 vccd1 vccd1 controller_627/HI la_data_out[9] sky130_fd_sc_hd__conb_1
Xcontroller_638 vssd1 vssd1 vccd1 vccd1 controller_638/HI la_data_out[20] sky130_fd_sc_hd__conb_1
XFILLER_0_28_261 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_28_283 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_1958_ _2002_/A vssd1 vssd1 vccd1 vccd1 _1958_/Y sky130_fd_sc_hd__inv_2
Xcontroller_649 vssd1 vssd1 vccd1 vccd1 controller_649/HI la_data_out[31] sky130_fd_sc_hd__conb_1
XFILLER_0_16_456 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_22_91 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_1889_ _2039_/A vssd1 vssd1 vccd1 vccd1 _1889_/Y sky130_fd_sc_hd__inv_2
XFILLER_0_16_489 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_31_459 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__1535__B1 _1541_/B1 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xinput117 data_in[58] vssd1 vssd1 vccd1 vccd1 _1515_/A1 sky130_fd_sc_hd__dlymetal6s2s_1
Xinput106 data_in[48] vssd1 vssd1 vccd1 vccd1 _1535_/A1 sky130_fd_sc_hd__buf_1
Xinput139 data_in[78] vssd1 vssd1 vccd1 vccd1 _1475_/A1 sky130_fd_sc_hd__buf_2
Xinput128 data_in[68] vssd1 vssd1 vccd1 vccd1 _1495_/A1 sky130_fd_sc_hd__buf_2
XPHY_112 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_101 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_39_537 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_47_570 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__2063__A _2069_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__1378__S hold26/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_50_713 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_34_253 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XANTENNA_hold972_A _2083_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_34_297 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_27_47 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_43_35 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XPHY_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_57_334 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_43_57 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_45_518 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__1288__S _1318_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_1812_ _2070_/Q _2248_/Q _2249_/Q vssd1 vssd1 vccd1 vccd1 _1812_/X sky130_fd_sc_hd__and3_1
X_1743_ _2181_/Q _1756_/B vssd1 vssd1 vccd1 vccd1 _1743_/X sky130_fd_sc_hd__and2_1
XFILLER_0_41_713 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_13_426 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_1674_ _2102_/Q _1677_/B vssd1 vssd1 vccd1 vccd1 _1674_/X sky130_fd_sc_hd__and2_1
Xhold316 hold316/A vssd1 vssd1 vccd1 vccd1 _1253_/B sky130_fd_sc_hd__dlygate4sd3_1
Xhold305 hold328/X vssd1 vssd1 vccd1 vccd1 hold305/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold349 _1487_/X vssd1 vssd1 vccd1 vccd1 hold349/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold338 hold356/X vssd1 vssd1 vccd1 vccd1 hold338/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold327 _1252_/X vssd1 vssd1 vccd1 vccd1 _2227_/D sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_40_256 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__1517__B1 _1529_/B1 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_21_470 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_610 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_632 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_621 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_643 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_676 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_665 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_654 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_698 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_687 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_2226_ _2239_/CLK _2226_/D _1966_/Y vssd1 vssd1 vccd1 vccd1 _2226_/Q sky130_fd_sc_hd__dfrtp_2
X_2157_ _2251_/CLK _2157_/D _1898_/Y vssd1 vssd1 vccd1 vccd1 _2157_/Q sky130_fd_sc_hd__dfrtp_1
XFILLER_0_16_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__1296__A2 _1529_/A2 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_2088_ _2168_/CLK _2088_/D _1831_/Y vssd1 vssd1 vccd1 vccd1 _2088_/Q sky130_fd_sc_hd__dfrtp_4
X_1108_ _2202_/Q _2110_/Q _1188_/S vssd1 vssd1 vccd1 vccd1 _1108_/X sky130_fd_sc_hd__mux2_1
XFILLER_0_48_312 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_1039_ hold571/X _1057_/A2 _1057_/B1 _1038_/X vssd1 vssd1 vccd1 vccd1 _2325_/D sky130_fd_sc_hd__a22o_1
XANTENNA_fanout606_A input262/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_44_573 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_44_562 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_16_286 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_31_234 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xhold872 _2271_/Q vssd1 vssd1 vccd1 vccd1 hold872/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold861 _2264_/Q vssd1 vssd1 vccd1 vccd1 hold861/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold850 _2280_/Q vssd1 vssd1 vccd1 vccd1 hold850/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold883 la_data_in[55] vssd1 vssd1 vccd1 vccd1 hold883/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold894 la_data_in[8] vssd1 vssd1 vccd1 vccd1 hold894/X sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA_clkbuf_leaf_16_wb_clk_i_A clkbuf_1_1__f_wb_clk_i/X vssd1 vssd1 vccd1 vccd1
+ sky130_fd_sc_hd__diode_2
XANTENNA__1287__A2 _1529_/A2 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__2058__A _2069_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_39_301 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__1897__A _2065_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_39_378 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_39_389 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_10_418 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_1390_ _1389_/X hold966/X _1435_/S vssd1 vssd1 vccd1 vccd1 _2181_/D sky130_fd_sc_hd__mux2_1
XFILLER_0_38_57 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_2011_ _2034_/A vssd1 vssd1 vccd1 vccd1 _2011_/Y sky130_fd_sc_hd__inv_2
XANTENNA__1278__A2 _1519_/A2 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_54_89 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_58_698 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_45_337 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_5_423 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_41_554 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xhold124 _1461_/X vssd1 vssd1 vccd1 vccd1 _2157_/D sky130_fd_sc_hd__dlygate4sd3_1
Xhold135 hold135/A vssd1 vssd1 vccd1 vccd1 _1343_/B sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA__1202__A2 _1202_/A2 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_13_245 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
Xhold113 hold79/X vssd1 vssd1 vccd1 vccd1 _1530_/S sky130_fd_sc_hd__buf_1
X_1726_ _2164_/Q _1766_/B vssd1 vssd1 vccd1 vccd1 _1726_/X sky130_fd_sc_hd__and2_1
Xhold102 _1613_/X vssd1 vssd1 vccd1 vccd1 hold102/X sky130_fd_sc_hd__dlygate4sd3_1
X_1657_ _2085_/Q _1680_/B vssd1 vssd1 vccd1 vccd1 _1657_/X sky130_fd_sc_hd__and2_1
Xhold146 hold146/A vssd1 vssd1 vccd1 vccd1 _1298_/B sky130_fd_sc_hd__dlygate4sd3_1
Xhold168 hold168/A vssd1 vssd1 vccd1 vccd1 _1208_/B sky130_fd_sc_hd__dlygate4sd3_1
Xhold157 _1609_/X vssd1 vssd1 vccd1 vccd1 hold157/X sky130_fd_sc_hd__dlygate4sd3_1
X_1588_ hold526/X hold981/X _1622_/S vssd1 vssd1 vccd1 vccd1 _2092_/D sky130_fd_sc_hd__mux2_1
Xfanout615 input262/X vssd1 vssd1 vccd1 vccd1 _2061_/A sky130_fd_sc_hd__clkbuf_8
Xfanout604 _1957_/A vssd1 vssd1 vccd1 vccd1 _1954_/A sky130_fd_sc_hd__buf_8
Xhold179 _1532_/X vssd1 vssd1 vccd1 vccd1 _2120_/D sky130_fd_sc_hd__dlygate4sd3_1
XTAP_440 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_451 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_473 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_462 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_484 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_495 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__1269__A2 _1519_/A2 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout556_A _1097_/B1 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_2209_ _2212_/CLK hold97/X _1949_/Y vssd1 vssd1 vccd1 vccd1 _2209_/Q sky130_fd_sc_hd__dfrtp_4
XFILLER_0_8_261 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_51_307 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_17_573 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_44_392 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_44_381 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_17_595 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_32_576 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
Xhold680 hold823/X vssd1 vssd1 vccd1 vccd1 hold680/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold691 hold862/X vssd1 vssd1 vccd1 vccd1 hold691/X sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA_hold935_A _2196_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_24_15 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_24_26 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_24_37 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_24_48 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_27_337 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XANTENNA_output475_A hold568/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_23_521 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_2_448 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_1511_ _1511_/A1 _1519_/A2 _1519_/B1 _2131_/Q hold500/X vssd1 vssd1 vccd1 vccd1 _1511_/X
+ sky130_fd_sc_hd__a221o_1
X_1442_ _1445_/A hold30/X vssd1 vssd1 vccd1 vccd1 hold31/A sky130_fd_sc_hd__and2_1
X_1373_ _1415_/A _1373_/B vssd1 vssd1 vccd1 vccd1 _1373_/X sky130_fd_sc_hd__and2_1
XANTENNA__1120__A1 _2104_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__1476__S _1504_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_26_370 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_26_392 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_14_587 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_1709_ _2137_/Q _1766_/B vssd1 vssd1 vccd1 vccd1 _1709_/X sky130_fd_sc_hd__and2_1
XTAP_281 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_270 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_292 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xclkbuf_leaf_5_wb_clk_i clkbuf_leaf_9_wb_clk_i/A vssd1 vssd1 vccd1 vccd1 _2182_/CLK
+ sky130_fd_sc_hd__clkbuf_16
XFILLER_0_49_495 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_36_167 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_36_189 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__1178__A1 _2075_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_32_373 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_32_384 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__1415__A _1415_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__1350__B2 _2195_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__1102__A1 _2113_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_35_69 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_51_46 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_1991_ _2008_/A vssd1 vssd1 vccd1 vccd1 _1991_/Y sky130_fd_sc_hd__inv_2
XFILLER_0_42_104 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_42_126 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_3_713 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_23_362 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_23_384 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_2_289 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_1425_ _1425_/A1 _1569_/A2 _1569_/B1 _2170_/Q hold117/X vssd1 vssd1 vccd1 vccd1 _1425_/X
+ sky130_fd_sc_hd__a221o_1
X_1356_ input15/X _1533_/A2 _1529_/B1 _2193_/Q hold276/X vssd1 vssd1 vccd1 vccd1 _1356_/X
+ sky130_fd_sc_hd__a221o_1
XANTENNA__1341__B2 _2198_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_1287_ input40/X _1529_/A2 _1529_/B1 _2216_/Q hold353/X vssd1 vssd1 vccd1 vccd1 _1287_/X
+ sky130_fd_sc_hd__a221o_1
XFILLER_0_46_421 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_18_123 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__1995__A _2002_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_46_465 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_14_340 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XANTENNA__1332__B2 _2201_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__2066__A _2069_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__1096__A0 _2208_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_49_292 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_24_159 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_20_365 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__1571__B2 _2101_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_2190_ _2194_/CLK _2190_/D _1930_/Y vssd1 vssd1 vccd1 vccd1 _2190_/Q sky130_fd_sc_hd__dfrtp_4
X_1210_ _1209_/X _2241_/Q _1252_/S vssd1 vssd1 vccd1 vccd1 _1210_/X sky130_fd_sc_hd__mux2_1
X_1141_ _2274_/Q _1189_/A2 _1189_/B1 _1140_/X vssd1 vssd1 vccd1 vccd1 _1141_/X sky130_fd_sc_hd__a22o_1
XANTENNA__1323__A1 input27/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__1323__B2 _2204_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_1072_ _2220_/Q hold994/X _1086_/S vssd1 vssd1 vccd1 vccd1 _1072_/X sky130_fd_sc_hd__mux2_1
XANTENNA__1087__B1 _1095_/B1 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_28_410 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_28_421 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_1974_ _1979_/A vssd1 vssd1 vccd1 vccd1 _1974_/Y sky130_fd_sc_hd__inv_2
XFILLER_0_7_337 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_7_359 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_16_638 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_43_468 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_11_310 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_23_192 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_24_693 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_30_129 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_46_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
Xhold17 hold17/A vssd1 vssd1 vccd1 vccd1 hold17/X sky130_fd_sc_hd__buf_1
Xhold28 hold28/A vssd1 vssd1 vccd1 vccd1 hold28/X sky130_fd_sc_hd__dlygate4sd3_1
X_1408_ _1407_/X hold953/X hold27/X vssd1 vssd1 vccd1 vccd1 _1408_/X sky130_fd_sc_hd__mux2_1
Xhold39 hold39/A vssd1 vssd1 vccd1 vccd1 hold39/X sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA__1314__B2 _2207_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_1339_ _1338_/X _2198_/Q _1372_/S vssd1 vssd1 vccd1 vccd1 _1339_/X sky130_fd_sc_hd__mux2_1
XANTENNA__1078__A0 _2217_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_46_251 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_46_284 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_34_402 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_34_413 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_15_671 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_30_641 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__1553__B2 _2110_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xoutput390 _1710_/X vssd1 vssd1 vccd1 vccd1 data_out[68] sky130_fd_sc_hd__buf_12
XANTENNA__1305__B2 _2210_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_16_16 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__1069__B1 _1097_/B1 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_37_251 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_4_307 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_37_262 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_52_265 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
Xhold509 hold773/X vssd1 vssd1 vccd1 vccd1 hold509/X sky130_fd_sc_hd__dlygate4sd3_1
X_1690_ _2118_/Q _1724_/B vssd1 vssd1 vccd1 vccd1 _1690_/X sky130_fd_sc_hd__and2_1
XFILLER_0_21_630 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_825 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_814 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_803 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_2311_ _2328_/CLK _2311_/D _2050_/Y vssd1 vssd1 vccd1 vccd1 _2311_/Q sky130_fd_sc_hd__dfrtp_1
XFILLER_0_20_173 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__1544__A1 _2114_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_858 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_847 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_836 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_20_195 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_869 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_2242_ _2322_/CLK _2242_/D _1982_/Y vssd1 vssd1 vccd1 vccd1 _2242_/Q sky130_fd_sc_hd__dfrtp_1
X_2173_ _2173_/CLK _2173_/D _1913_/Y vssd1 vssd1 vccd1 vccd1 _2173_/Q sky130_fd_sc_hd__dfrtp_4
X_1124_ _2194_/Q _2102_/Q _1156_/S vssd1 vssd1 vccd1 vccd1 _1124_/X sky130_fd_sc_hd__mux2_1
X_1055_ hold590/X _1095_/A2 _1057_/B1 _1054_/X vssd1 vssd1 vccd1 vccd1 _2317_/D sky130_fd_sc_hd__a22o_1
XFILLER_0_18_7 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_28_240 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xcontroller_628 vssd1 vssd1 vccd1 vccd1 controller_628/HI la_data_out[10] sky130_fd_sc_hd__conb_1
Xcontroller_639 vssd1 vssd1 vccd1 vccd1 controller_639/HI la_data_out[21] sky130_fd_sc_hd__conb_1
XFILLER_0_16_413 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_1957_ _1957_/A vssd1 vssd1 vccd1 vccd1 _1957_/Y sky130_fd_sc_hd__inv_2
XFILLER_0_16_468 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_28_295 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_1888_ _2039_/A vssd1 vssd1 vccd1 vccd1 _1888_/Y sky130_fd_sc_hd__inv_2
XFILLER_0_43_287 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_43_254 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_31_449 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__1484__S _1504_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__1535__A1 _1535_/A1 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__1535__B2 _2119_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xinput118 data_in[59] vssd1 vssd1 vccd1 vccd1 _1513_/A1 sky130_fd_sc_hd__buf_1
Xinput107 data_in[49] vssd1 vssd1 vccd1 vccd1 _1533_/A1 sky130_fd_sc_hd__buf_1
XANTENNA_fanout586_A _1112_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xinput129 data_in[69] vssd1 vssd1 vccd1 vccd1 _1493_/A1 sky130_fd_sc_hd__clkbuf_2
XANTENNA__1299__B1 _1529_/B1 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_39_505 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XPHY_113 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_102 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__1471__B1 _1541_/B1 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_35_700 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_34_265 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_34_287 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA_hold965_A _2073_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__1526__A1 _2123_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_27_15 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_57_302 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_43_69 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XPHY_4 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_45_508 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_1811_ _1811_/A _1811_/B vssd1 vssd1 vccd1 vccd1 _2156_/D sky130_fd_sc_hd__nor2_1
XFILLER_0_38_571 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_4_104 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_1742_ _2180_/Q _1756_/B vssd1 vssd1 vccd1 vccd1 _1742_/X sky130_fd_sc_hd__and2_1
XFILLER_0_13_405 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_1673_ _2101_/Q _1677_/B vssd1 vssd1 vccd1 vccd1 _1673_/X sky130_fd_sc_hd__and2_1
Xhold306 hold306/A vssd1 vssd1 vccd1 vccd1 _1259_/B sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_13_438 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_13_449 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xhold317 _1253_/X vssd1 vssd1 vccd1 vccd1 hold317/X sky130_fd_sc_hd__buf_1
Xhold328 la_data_in[62] vssd1 vssd1 vccd1 vccd1 hold328/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold339 hold339/A vssd1 vssd1 vccd1 vccd1 _1274_/B sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA__1517__A1 _1517_/A1 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_21_482 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_600 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_0_365 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_611 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_633 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_622 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_677 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_666 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_655 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_644 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_699 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_688 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_2225_ _2225_/CLK _2225_/D _1965_/Y vssd1 vssd1 vccd1 vccd1 _2225_/Q sky130_fd_sc_hd__dfrtp_2
X_2156_ _2156_/D _1813_/X vssd1 vssd1 vccd1 vccd1 _2156_/Q sky130_fd_sc_hd__dlxtn_1
X_2087_ _2168_/CLK _2087_/D _1830_/Y vssd1 vssd1 vccd1 vccd1 _2087_/Q sky130_fd_sc_hd__dfrtp_4
X_1107_ hold763/X _1139_/A2 _1139_/B1 _1106_/X vssd1 vssd1 vccd1 vccd1 _2291_/D sky130_fd_sc_hd__a22o_1
X_1038_ _2237_/Q _2145_/Q _1038_/S vssd1 vssd1 vccd1 vccd1 _1038_/X sky130_fd_sc_hd__mux2_2
XFILLER_0_36_519 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_8_432 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_44_585 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_16_298 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
Xhold851 _2324_/Q vssd1 vssd1 vccd1 vccd1 hold851/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold873 la_data_in[9] vssd1 vssd1 vccd1 vccd1 hold873/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold840 la_data_in[0] vssd1 vssd1 vccd1 vccd1 hold840/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold862 _2257_/Q vssd1 vssd1 vccd1 vccd1 hold862/X sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_31_279 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xhold884 _1282_/X vssd1 vssd1 vccd1 vccd1 _2217_/D sky130_fd_sc_hd__dlygate4sd3_1
Xhold895 _1423_/X vssd1 vssd1 vccd1 vccd1 _2170_/D sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_54_305 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_50_533 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_50_511 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA_clkbuf_leaf_1_wb_clk_i_A clkbuf_leaf_9_wb_clk_i/A vssd1 vssd1 vccd1 vccd1
+ sky130_fd_sc_hd__diode_2
XFILLER_0_22_268 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_38_69 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__1380__C1 hold525/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_2010_ _2033_/A vssd1 vssd1 vccd1 vccd1 _2010_/Y sky130_fd_sc_hd__inv_2
XFILLER_0_57_110 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_18_508 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_45_349 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_26_530 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_5_446 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_53_371 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_1725_ _2163_/Q _1725_/B vssd1 vssd1 vccd1 vccd1 _1725_/X sky130_fd_sc_hd__and2_2
Xhold125 hold193/X vssd1 vssd1 vccd1 vccd1 hold125/X sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_13_257 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
Xhold103 _1614_/X vssd1 vssd1 vccd1 vccd1 _2079_/D sky130_fd_sc_hd__dlygate4sd3_1
Xhold114 _1542_/X vssd1 vssd1 vccd1 vccd1 _2115_/D sky130_fd_sc_hd__dlygate4sd3_1
Xhold147 _1298_/X vssd1 vssd1 vccd1 vccd1 hold147/X sky130_fd_sc_hd__buf_1
Xhold158 _1610_/X vssd1 vssd1 vccd1 vccd1 _2081_/D sky130_fd_sc_hd__dlygate4sd3_1
Xhold136 _1343_/X vssd1 vssd1 vccd1 vccd1 hold136/X sky130_fd_sc_hd__dlymetal6s2s_1
X_1656_ _2084_/Q _1680_/B vssd1 vssd1 vccd1 vccd1 _1656_/X sky130_fd_sc_hd__and2_1
X_1587_ input78/X _1619_/A2 _1619_/B1 _2093_/Q hold525/X vssd1 vssd1 vccd1 vccd1 _1587_/X
+ sky130_fd_sc_hd__a221o_1
Xhold169 _1208_/X vssd1 vssd1 vccd1 vccd1 hold169/X sky130_fd_sc_hd__buf_1
Xfanout605 _1949_/A vssd1 vssd1 vccd1 vccd1 _1957_/A sky130_fd_sc_hd__buf_4
XTAP_430 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_441 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xfanout616 _2039_/A vssd1 vssd1 vccd1 vccd1 _1979_/A sky130_fd_sc_hd__buf_8
XANTENNA__1371__C1 hold208/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_452 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_474 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_463 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_485 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_496 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_2208_ _2269_/CLK hold61/X _1948_/Y vssd1 vssd1 vccd1 vccd1 _2208_/Q sky130_fd_sc_hd__dfrtp_4
X_2139_ _2239_/CLK _2139_/D _1882_/Y vssd1 vssd1 vccd1 vccd1 _2139_/Q sky130_fd_sc_hd__dfrtp_1
XFILLER_0_8_273 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA_hold127_A _1373_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_8_295 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_17_552 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_32_599 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_12_290 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
Xhold670 hold866/X vssd1 vssd1 vccd1 vccd1 hold670/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold681 hold812/X vssd1 vssd1 vccd1 vccd1 hold681/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold692 hold822/X vssd1 vssd1 vccd1 vccd1 hold692/X sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA__1362__C1 hold223/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__2069__A _2069_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_59_419 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_39_121 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_55_614 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_27_316 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_27_349 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_2_405 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_23_511 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_23_544 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_1510_ _1509_/X hold914/X _1520_/S vssd1 vssd1 vccd1 vccd1 _2131_/D sky130_fd_sc_hd__mux2_1
XFILLER_0_50_363 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_49_68 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_49_57 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_1441_ _1440_/X _2164_/Q hold27/X vssd1 vssd1 vccd1 vccd1 hold28/A sky130_fd_sc_hd__mux2_1
XANTENNA__1353__C1 hold244/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_1372_ _1371_/X _2187_/Q _1372_/S vssd1 vssd1 vccd1 vccd1 _1372_/X sky130_fd_sc_hd__mux2_1
XFILLER_0_58_474 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_18_305 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_45_124 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_45_113 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_18_327 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_14_533 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__1187__A2 _1189_/A2 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_41_385 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_1708_ _2136_/Q _1766_/B vssd1 vssd1 vccd1 vccd1 _1708_/X sky130_fd_sc_hd__and2_1
XFILLER_0_41_396 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_1639_ _1445_/A _2155_/D _1638_/X vssd1 vssd1 vccd1 vccd1 _2248_/D sky130_fd_sc_hd__o21a_1
XANTENNA__1492__S _1520_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__1344__C1 hold136/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_260 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_282 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_271 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_293 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_hold244_A _1352_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_49_463 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_9_593 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_51_116 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_17_393 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_20_503 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_20_536 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_20_547 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__1583__C1 hold127/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_35_15 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_1990_ _2008_/A vssd1 vssd1 vccd1 vccd1 _1990_/Y sky130_fd_sc_hd__inv_2
XFILLER_0_7_508 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_27_113 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_28_636 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_27_157 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_43_628 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_15_319 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_42_138 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__1169__A2 _1183_/A2 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_50_182 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_11_558 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_1424_ _1445_/A _1424_/B vssd1 vssd1 vccd1 vccd1 _1424_/X sky130_fd_sc_hd__and2_1
X_1355_ _1415_/A _1355_/B vssd1 vssd1 vccd1 vccd1 _1355_/X sky130_fd_sc_hd__and2_1
X_1286_ _1310_/A _1286_/B vssd1 vssd1 vccd1 vccd1 _1286_/X sky130_fd_sc_hd__and2_1
XFILLER_0_25_81 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_19_625 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_46_433 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_46_411 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_46_477 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_6_530 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_6_585 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_14_352 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__1565__C1 hold106/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__1332__A2 _1197_/D vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_37_411 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_25_617 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_25_628 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__1571__A2 _1623_/A2 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__1323__A2 _1197_/D vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_1140_ _2186_/Q _2094_/Q _1178_/S vssd1 vssd1 vccd1 vccd1 _1140_/X sky130_fd_sc_hd__mux2_1
X_1071_ hold575/X _1097_/A2 _1097_/B1 _1070_/X vssd1 vssd1 vccd1 vccd1 _2309_/D sky130_fd_sc_hd__a22o_1
XFILLER_0_47_208 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_1973_ _1979_/A vssd1 vssd1 vccd1 vccd1 _1973_/Y sky130_fd_sc_hd__inv_2
XFILLER_0_28_455 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_7_349 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__1100__S _1188_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_28_477 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_31_609 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_11_333 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xhold29 la_data_in[1] vssd1 vssd1 vccd1 vccd1 hold29/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold18 hold18/A vssd1 vssd1 vccd1 vccd1 hold18/X sky130_fd_sc_hd__dlygate4sd3_1
X_1407_ _1407_/A1 _1003_/Y _1569_/B1 _2176_/Q hold219/X vssd1 vssd1 vccd1 vccd1 _1407_/X
+ sky130_fd_sc_hd__a221o_1
XANTENNA__1314__A2 _1197_/D vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_39_3 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_1338_ input21/X _1533_/A2 _1533_/B1 _2199_/Q hold344/X vssd1 vssd1 vccd1 vccd1 _1338_/X
+ sky130_fd_sc_hd__a221o_1
X_1269_ input47/X _1519_/A2 _1519_/B1 _2222_/Q hold463/X vssd1 vssd1 vccd1 vccd1 _1269_/X
+ sky130_fd_sc_hd__a221o_1
XANTENNA__1078__A1 _2125_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout531_A _1097_/A2 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_19_422 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_46_241 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_19_466 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_46_296 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_6_360 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
Xoutput380 _1701_/X vssd1 vssd1 vccd1 vccd1 data_out[59] sky130_fd_sc_hd__buf_12
XANTENNA__1553__A2 _1637_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xoutput391 _1711_/X vssd1 vssd1 vccd1 vccd1 data_out[69] sky130_fd_sc_hd__buf_12
XANTENNA__1305__A2 _1527_/A2 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_29_219 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_52_233 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_4_319 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_52_277 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_40_406 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_20_141 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_21_642 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_826 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_815 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_804 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_2310_ _2315_/CLK _2310_/D _2049_/Y vssd1 vssd1 vccd1 vccd1 _2310_/Q sky130_fd_sc_hd__dfrtp_1
XTAP_859 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_848 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_837 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_2241_ _2322_/CLK _2241_/D _1981_/Y vssd1 vssd1 vccd1 vccd1 _2241_/Q sky130_fd_sc_hd__dfrtp_1
X_2172_ _2173_/CLK _2172_/D _1912_/Y vssd1 vssd1 vccd1 vccd1 _2172_/Q sky130_fd_sc_hd__dfrtp_4
X_1123_ hold647/X _1183_/A2 _1183_/B1 _1122_/X vssd1 vssd1 vccd1 vccd1 _2283_/D sky130_fd_sc_hd__a22o_1
X_1054_ _2229_/Q _2137_/Q _1094_/S vssd1 vssd1 vccd1 vccd1 _1054_/X sky130_fd_sc_hd__mux2_1
XFILLER_0_7_102 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_1956_ _1957_/A vssd1 vssd1 vccd1 vccd1 _1956_/Y sky130_fd_sc_hd__inv_2
Xcontroller_618 vssd1 vssd1 vccd1 vccd1 controller_618/HI la_data_out[0] sky130_fd_sc_hd__conb_1
Xcontroller_629 vssd1 vssd1 vccd1 vccd1 controller_629/HI la_data_out[11] sky130_fd_sc_hd__conb_1
X_1887_ _1979_/A vssd1 vssd1 vccd1 vccd1 _1887_/Y sky130_fd_sc_hd__inv_2
XFILLER_0_24_480 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__1535__A2 _1197_/D vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xinput108 data_in[4] vssd1 vssd1 vccd1 vccd1 _1623_/A1 sky130_fd_sc_hd__buf_1
Xinput119 data_in[5] vssd1 vssd1 vccd1 vccd1 _1621_/A1 sky130_fd_sc_hd__clkbuf_1
XANTENNA_fanout579_A _1527_/B1 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__1299__B2 _2212_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XPHY_114 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_103 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__1471__A1 _1471_/A1 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__1471__B2 _2151_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_47_561 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_35_712 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_34_222 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_15_491 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_22_439 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA_hold958_A _2075_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_43_15 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XPHY_5 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__1462__A1 _1527_/A2 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_1810_ _1810_/A _1810_/B _1810_/C _1810_/D vssd1 vssd1 vccd1 vccd1 _1811_/B sky130_fd_sc_hd__or4_1
XFILLER_0_26_701 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_38_561 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_38_583 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_1741_ _2179_/Q _1756_/B vssd1 vssd1 vccd1 vccd1 _1741_/X sky130_fd_sc_hd__and2_1
X_1672_ _2100_/Q _1677_/B vssd1 vssd1 vccd1 vccd1 _1672_/X sky130_fd_sc_hd__and2_1
Xhold307 _1259_/X vssd1 vssd1 vccd1 vccd1 hold307/X sky130_fd_sc_hd__buf_1
XFILLER_0_40_203 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
Xhold329 _1261_/X vssd1 vssd1 vccd1 vccd1 _2224_/D sky130_fd_sc_hd__dlygate4sd3_1
Xhold318 _1254_/X vssd1 vssd1 vccd1 vccd1 hold318/X sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA__1517__A2 _1529_/A2 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_21_461 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_601 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_612 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_634 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_623 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_667 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_656 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_645 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_2224_ _2224_/CLK _2224_/D _1964_/Y vssd1 vssd1 vccd1 vccd1 _2224_/Q sky130_fd_sc_hd__dfrtp_2
XTAP_689 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_678 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_2155_ _2155_/D _1445_/A vssd1 vssd1 vccd1 vccd1 _2155_/Q sky130_fd_sc_hd__dlxtn_1
XANTENNA__1150__A0 _2181_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_17_60 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_1106_ hold976/X _2111_/Q _1188_/S vssd1 vssd1 vccd1 vccd1 _1106_/X sky130_fd_sc_hd__mux2_1
X_2086_ _2168_/CLK _2086_/D _1829_/Y vssd1 vssd1 vccd1 vccd1 _2086_/Q sky130_fd_sc_hd__dfrtp_4
X_1037_ hold637/X _1095_/A2 _1095_/B1 _1036_/X vssd1 vssd1 vccd1 vccd1 _2326_/D sky130_fd_sc_hd__a22o_1
XFILLER_0_16_200 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_44_542 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_44_531 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_44_553 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_1939_ _1954_/A vssd1 vssd1 vccd1 vccd1 _1939_/Y sky130_fd_sc_hd__inv_2
Xinput90 data_in[33] vssd1 vssd1 vccd1 vccd1 input90/X sky130_fd_sc_hd__clkbuf_1
Xhold830 _2260_/Q vssd1 vssd1 vccd1 vccd1 hold830/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold863 _2308_/Q vssd1 vssd1 vccd1 vccd1 hold863/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold852 _2319_/Q vssd1 vssd1 vccd1 vccd1 hold852/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold841 _1447_/X vssd1 vssd1 vccd1 vccd1 _2162_/D sky130_fd_sc_hd__dlygate4sd3_1
Xhold885 _2327_/Q vssd1 vssd1 vccd1 vccd1 hold885/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold896 _2325_/Q vssd1 vssd1 vccd1 vccd1 hold896/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold874 _1420_/X vssd1 vssd1 vccd1 vccd1 _2171_/D sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA__1141__B1 _1189_/B1 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__1444__A1 _2163_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_27_509 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_54_328 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_35_575 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_22_214 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_50_589 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_50_578 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_38_15 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XANTENNA__1380__B1 _1529_/B1 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_54_25 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__1132__A0 _2190_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_54_69 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__1435__A1 hold979/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_45_317 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_26_553 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_13_225 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_1724_ _2162_/Q _1724_/B vssd1 vssd1 vccd1 vccd1 _1724_/X sky130_fd_sc_hd__and2_2
Xhold126 hold126/A vssd1 vssd1 vccd1 vccd1 _1373_/B sky130_fd_sc_hd__dlygate4sd3_1
Xhold104 hold144/X vssd1 vssd1 vccd1 vccd1 hold104/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold115 hold149/X vssd1 vssd1 vccd1 vccd1 hold115/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold137 _1563_/X vssd1 vssd1 vccd1 vccd1 hold137/X sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_41_578 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xhold159 hold844/X vssd1 vssd1 vccd1 vccd1 hold42/A sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_13_269 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xhold148 _1533_/X vssd1 vssd1 vccd1 vccd1 hold148/X sky130_fd_sc_hd__dlygate4sd3_1
X_1655_ _2083_/Q _1725_/B vssd1 vssd1 vccd1 vccd1 _1655_/X sky130_fd_sc_hd__and2_1
XFILLER_0_0_141 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xfanout606 input262/X vssd1 vssd1 vccd1 vccd1 _1949_/A sky130_fd_sc_hd__buf_8
X_1586_ _1585_/X hold990/X _1632_/S vssd1 vssd1 vccd1 vccd1 _2093_/D sky130_fd_sc_hd__mux2_1
XTAP_420 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_431 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_442 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xfanout617 input262/X vssd1 vssd1 vccd1 vccd1 _2039_/A sky130_fd_sc_hd__clkbuf_8
XTAP_453 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_475 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_464 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_2207_ _2269_/CLK hold14/X _1947_/Y vssd1 vssd1 vccd1 vccd1 _2207_/Q sky130_fd_sc_hd__dfrtp_4
XTAP_486 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_497 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_21_3 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XANTENNA__1123__B1 _1183_/B1 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_2138_ _2239_/CLK _2138_/D _1881_/Y vssd1 vssd1 vccd1 vccd1 _2138_/Q sky130_fd_sc_hd__dfrtp_1
X_2069_ _2069_/A vssd1 vssd1 vccd1 vccd1 _2069_/Y sky130_fd_sc_hd__inv_2
XFILLER_0_48_133 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA_fanout611_A input262/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_17_564 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_32_589 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xhold660 hold802/X vssd1 vssd1 vccd1 vccd1 hold660/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold671 hold834/X vssd1 vssd1 vccd1 vccd1 hold671/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold682 hold798/X vssd1 vssd1 vccd1 vccd1 hold682/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold693 hold813/X vssd1 vssd1 vccd1 vccd1 hold693/X sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA__1114__A0 _2199_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__1701__B _1715_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__1417__A1 _2172_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_39_133 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_27_306 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_27_328 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_54_169 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_54_158 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_54_147 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_35_361 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_23_556 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_50_397 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_1440_ _1440_/A1 _1637_/B _1545_/B1 _2165_/Q hold17/X vssd1 vssd1 vccd1 vccd1 _1440_/X
+ sky130_fd_sc_hd__a221o_1
X_1371_ input9/X _1533_/A2 _1533_/B1 _2188_/Q hold208/X vssd1 vssd1 vccd1 vccd1 _1371_/X
+ sky130_fd_sc_hd__a221o_1
XANTENNA__1353__B1 _1529_/B1 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_4_38 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_46_626 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_18_339 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_45_169 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_45_147 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_26_361 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_53_191 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_30_82 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_1707_ _2135_/Q _1761_/B vssd1 vssd1 vccd1 vccd1 _1707_/X sky130_fd_sc_hd__and2_1
XFILLER_0_41_353 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_1638_ _2248_/Q _2249_/Q _2161_/Q vssd1 vssd1 vccd1 vccd1 _1638_/X sky130_fd_sc_hd__or3_1
X_1569_ input88/X _1569_/A2 _1569_/B1 _2102_/Q hold244/X vssd1 vssd1 vccd1 vccd1 _1569_/X
+ sky130_fd_sc_hd__a221o_1
XTAP_250 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_39_80 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_283 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_272 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_261 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_294 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_fanout561_A _1569_/A2 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_49_475 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_37_615 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_37_626 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_36_136 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_32_353 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__1583__B1 _1623_/B1 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xhold490 la_data_in[83] vssd1 vssd1 vccd1 vccd1 hold490/X sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA_hold940_A _2104_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_27_103 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_27_169 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA_output480_A hold647/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_23_353 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_23_375 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_50_194 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_1423_ _1422_/X _2170_/Q hold27/X vssd1 vssd1 vccd1 vccd1 _1423_/X sky130_fd_sc_hd__mux2_1
XANTENNA__1326__B1 _1541_/B1 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_1354_ _1353_/X hold941/X _1372_/S vssd1 vssd1 vccd1 vccd1 _2193_/D sky130_fd_sc_hd__mux2_1
X_1285_ _1284_/X _2216_/Q _1318_/S vssd1 vssd1 vccd1 vccd1 _1285_/X sky130_fd_sc_hd__mux2_1
Xclkbuf_leaf_13_wb_clk_i clkbuf_1_1__f_wb_clk_i/X vssd1 vssd1 vccd1 vccd1 _2238_/CLK
+ sky130_fd_sc_hd__clkbuf_16
XANTENNA__1629__B2 _2072_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_19_604 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_58_283 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_18_103 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_19_637 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_19_648 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_46_456 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_46_445 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_27_670 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_26_191 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA_clkbuf_leaf_25_wb_clk_i_A clkbuf_leaf_9_wb_clk_i/A vssd1 vssd1 vccd1 vccd1
+ sky130_fd_sc_hd__diode_2
XANTENNA__1565__B1 _1569_/B1 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__1317__B1 _1541_/B1 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_52_404 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_9_391 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA_hold988_A _2172_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_32_150 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_33_651 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_20_345 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_20_356 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_32_194 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__1308__B1 _1541_/B1 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_1070_ _2221_/Q _2129_/Q _1086_/S vssd1 vssd1 vccd1 vccd1 _1070_/X sky130_fd_sc_hd__mux2_1
XANTENNA__1087__A2 _1095_/A2 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_7_306 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_1972_ _1979_/A vssd1 vssd1 vccd1 vccd1 _1972_/Y sky130_fd_sc_hd__inv_2
XFILLER_0_43_426 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_16_629 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_28_489 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_43_437 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_24_662 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_23_161 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_1406_ _1415_/A _1406_/B vssd1 vssd1 vccd1 vccd1 _1406_/X sky130_fd_sc_hd__and2_1
Xhold19 hold19/A vssd1 vssd1 vccd1 vccd1 hold19/X sky130_fd_sc_hd__dlygate4sd3_1
X_1337_ _1349_/A _1337_/B vssd1 vssd1 vccd1 vccd1 _1337_/X sky130_fd_sc_hd__and2_1
XANTENNA__1352__A _1415_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_1268_ _1271_/A _1268_/B vssd1 vssd1 vccd1 vccd1 _1268_/X sky130_fd_sc_hd__and2_1
X_1199_ hold2/X _1198_/X _1197_/X vssd1 vssd1 vccd1 vccd1 hold3/A sky130_fd_sc_hd__a21bo_1
XANTENNA__1483__C1 hold443/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_38_209 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__1498__S _1504_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout524_A hold26/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_46_253 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_19_489 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_15_662 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_21_109 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_42_470 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_14_183 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_30_621 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
Xoutput370 _1646_/X vssd1 vssd1 vccd1 vccd1 data_out[4] sky130_fd_sc_hd__buf_12
Xoutput381 _1647_/X vssd1 vssd1 vccd1 vccd1 data_out[5] sky130_fd_sc_hd__buf_12
Xoutput392 _1648_/X vssd1 vssd1 vccd1 vccd1 data_out[6] sky130_fd_sc_hd__buf_12
XANTENNA__1069__A2 _1097_/A2 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_37_275 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_40_418 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_52_289 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_21_621 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__1529__B1 _1529_/B1 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_20_120 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_21_665 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_816 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_805 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_0_559 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_20_153 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_849 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_57_47 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_838 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_827 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_20_197 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_2240_ _2322_/CLK _2240_/D _1980_/Y vssd1 vssd1 vccd1 vccd1 _2240_/Q sky130_fd_sc_hd__dfrtp_1
X_2171_ _2173_/CLK _2171_/D _1911_/Y vssd1 vssd1 vccd1 vccd1 _2171_/Q sky130_fd_sc_hd__dfrtp_4
X_1122_ _2195_/Q _2103_/Q _1178_/S vssd1 vssd1 vccd1 vccd1 _1122_/X sky130_fd_sc_hd__mux2_1
X_1053_ hold591/X _1057_/A2 _1057_/B1 _1052_/X vssd1 vssd1 vccd1 vccd1 _2318_/D sky130_fd_sc_hd__a22o_1
XANTENNA__1900__A _1913_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_1955_ _1957_/A vssd1 vssd1 vccd1 vccd1 _1955_/Y sky130_fd_sc_hd__inv_2
Xcontroller_619 vssd1 vssd1 vccd1 vccd1 controller_619/HI la_data_out[1] sky130_fd_sc_hd__conb_1
XFILLER_0_16_404 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_28_253 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_22_94 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_28_286 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_1886_ _1979_/A vssd1 vssd1 vccd1 vccd1 _1886_/Y sky130_fd_sc_hd__inv_2
XFILLER_0_43_278 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
Xinput109 data_in[50] vssd1 vssd1 vccd1 vccd1 _1531_/A1 sky130_fd_sc_hd__buf_1
XFILLER_0_51_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__1299__A2 _1529_/A2 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_2_93 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XPHY_115 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_104 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_47_551 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_19_220 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__1471__A2 _1197_/D vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_15_481 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_34_278 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_30_473 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_30_495 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__1704__B _1715_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_43_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XPHY_6 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_57_337 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_26_713 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_25_234 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_1740_ _2178_/Q _1761_/B vssd1 vssd1 vccd1 vccd1 _1740_/X sky130_fd_sc_hd__and2_1
X_1671_ _2099_/Q _1677_/B vssd1 vssd1 vccd1 vccd1 _1671_/X sky130_fd_sc_hd__and2_1
Xhold308 _1507_/X vssd1 vssd1 vccd1 vccd1 hold308/X sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_40_215 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
Xhold319 la_data_in[51] vssd1 vssd1 vccd1 vccd1 hold319/X sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_40_259 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_602 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_613 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_624 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_668 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_657 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_635 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_646 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_2223_ _2223_/CLK _2223_/D _1963_/Y vssd1 vssd1 vccd1 vccd1 _2223_/Q sky130_fd_sc_hd__dfrtp_4
XTAP_679 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__1106__S _1188_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_2154_ _2328_/CLK _2154_/D _1897_/Y vssd1 vssd1 vccd1 vccd1 _2154_/Q sky130_fd_sc_hd__dfrtp_1
XANTENNA__1150__A1 _2089_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_1105_ hold620/X _1139_/A2 _1139_/B1 _1104_/X vssd1 vssd1 vccd1 vccd1 _2292_/D sky130_fd_sc_hd__a22o_1
X_2085_ _2106_/CLK _2085_/D _1828_/Y vssd1 vssd1 vccd1 vccd1 _2085_/Q sky130_fd_sc_hd__dfrtp_4
X_1036_ _2238_/Q _2146_/Q _1086_/S vssd1 vssd1 vccd1 vccd1 _1036_/X sky130_fd_sc_hd__mux2_1
XFILLER_0_17_713 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_44_576 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_44_565 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_16_256 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_1938_ _1954_/A vssd1 vssd1 vccd1 vccd1 _1938_/Y sky130_fd_sc_hd__inv_2
X_1869_ _2002_/A vssd1 vssd1 vccd1 vccd1 _1869_/Y sky130_fd_sc_hd__inv_2
Xinput91 data_in[34] vssd1 vssd1 vccd1 vccd1 input91/X sky130_fd_sc_hd__clkbuf_1
Xinput80 data_in[24] vssd1 vssd1 vccd1 vccd1 input80/X sky130_fd_sc_hd__buf_1
Xhold820 _2282_/Q vssd1 vssd1 vccd1 vccd1 hold820/X sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_31_237 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
Xhold842 la_data_in[12] vssd1 vssd1 vccd1 vccd1 hold842/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold853 _2321_/Q vssd1 vssd1 vccd1 vccd1 hold853/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold864 _2259_/Q vssd1 vssd1 vccd1 vccd1 hold864/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold831 _2283_/Q vssd1 vssd1 vccd1 vccd1 hold831/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold886 la_data_in[39] vssd1 vssd1 vccd1 vccd1 hold886/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold875 _2304_/Q vssd1 vssd1 vccd1 vccd1 hold875/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold897 _2289_/Q vssd1 vssd1 vccd1 vccd1 hold897/X sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_39_304 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_39_315 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_39_337 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_47_381 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__1601__C1 hold132/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_35_587 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XANTENNA_hold970_A _2180_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_38_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__1380__B2 _2185_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_54_15 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__1132__A1 _2098_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_output406_A _1724_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_45_329 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_5_426 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_53_362 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_41_513 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_41_502 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_1723_ _2151_/Q _1766_/B vssd1 vssd1 vccd1 vccd1 _1723_/X sky130_fd_sc_hd__and2_2
XFILLER_0_41_557 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xhold105 hold105/A vssd1 vssd1 vccd1 vccd1 _1346_/B sky130_fd_sc_hd__dlygate4sd3_1
Xhold116 hold116/A vssd1 vssd1 vccd1 vccd1 _1424_/B sky130_fd_sc_hd__dlygate4sd3_1
Xhold149 hold917/X vssd1 vssd1 vccd1 vccd1 hold149/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold138 la_data_in[15] vssd1 vssd1 vccd1 vccd1 hold138/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold127 _1373_/X vssd1 vssd1 vccd1 vccd1 hold127/X sky130_fd_sc_hd__dlymetal6s2s_1
X_1654_ _2082_/Q _1725_/B vssd1 vssd1 vccd1 vccd1 _1654_/X sky130_fd_sc_hd__and2_1
XFILLER_0_21_281 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_1585_ input79/X _1623_/A2 _1623_/B1 _2094_/Q hold536/X vssd1 vssd1 vccd1 vccd1 _1585_/X
+ sky130_fd_sc_hd__a221o_1
Xfanout607 _2034_/A vssd1 vssd1 vccd1 vccd1 _2008_/A sky130_fd_sc_hd__buf_8
XTAP_410 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_421 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_432 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__1371__B2 _2188_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_443 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_454 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_476 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_465 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_2206_ _2212_/CLK _2206_/D _1946_/Y vssd1 vssd1 vccd1 vccd1 _2206_/Q sky130_fd_sc_hd__dfrtp_4
XFILLER_0_28_71 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_28_82 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_487 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_498 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__1123__A1 hold647/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_14_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_2137_ _2322_/CLK _2137_/D _1880_/Y vssd1 vssd1 vccd1 vccd1 _2137_/Q sky130_fd_sc_hd__dfrtp_1
X_2068_ _2069_/A vssd1 vssd1 vccd1 vccd1 _2068_/Y sky130_fd_sc_hd__inv_2
X_1019_ _1455_/A hold561/X hold778/X _1017_/X _0974_/X vssd1 vssd1 vccd1 vccd1 _1204_/B
+ sky130_fd_sc_hd__a32o_1
XFILLER_0_48_189 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA_fanout604_A _1957_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_17_576 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_32_557 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
Xhold661 hold876/X vssd1 vssd1 vccd1 vccd1 hold661/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold650 hold699/X vssd1 vssd1 vccd1 vccd1 hold650/X sky130_fd_sc_hd__clkbuf_2
Xhold672 hold811/X vssd1 vssd1 vccd1 vccd1 hold672/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold694 hold864/X vssd1 vssd1 vccd1 vccd1 hold694/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold683 hold801/X vssd1 vssd1 vccd1 vccd1 hold683/X sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA__1362__B2 _2191_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__1114__A1 _2107_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_39_101 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_39_145 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_39_167 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_54_137 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_35_373 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_2_418 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_50_365 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_49_15 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_1370_ _1415_/A _1370_/B vssd1 vssd1 vccd1 vccd1 _1370_/X sky130_fd_sc_hd__and2_1
XANTENNA__1353__B2 _2194_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_18_318 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_45_159 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_6_713 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_26_373 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_53_181 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_5_278 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_26_395 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA_clkbuf_leaf_15_wb_clk_i_A clkbuf_1_1__f_wb_clk_i/X vssd1 vssd1 vccd1 vccd1
+ sky130_fd_sc_hd__diode_2
X_1706_ _2134_/Q _1715_/B vssd1 vssd1 vccd1 vccd1 _1706_/X sky130_fd_sc_hd__and2_1
X_1637_ _1637_/A _1637_/B vssd1 vssd1 vccd1 vccd1 _2155_/D sky130_fd_sc_hd__nor2_1
XANTENNA__1355__A _1415_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_1568_ hold407/X hold921/X hold81/X vssd1 vssd1 vccd1 vccd1 _2102_/D sky130_fd_sc_hd__mux2_1
XANTENNA__1344__B2 _2197_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_251 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_240 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_284 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_273 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_262 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_1499_ _1499_/A1 _1463_/B _1499_/B1 _2137_/Q hold312/X vssd1 vssd1 vccd1 vccd1 _1499_/X
+ sky130_fd_sc_hd__a221o_1
XTAP_295 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_55_80 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA_fanout554_A _1157_/B1 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_49_498 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_36_104 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_44_192 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_32_365 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_32_387 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__1583__B2 _2095_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xhold480 la_data_in[76] vssd1 vssd1 vccd1 vccd1 hold480/X sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_3_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xhold491 hold491/A vssd1 vssd1 vccd1 vccd1 _0977_/B sky130_fd_sc_hd__dlymetal6s2s_1
XANTENNA__1335__B2 _2200_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_hold933_A _2103_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__1099__B1 _1157_/B1 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_59_207 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_55_446 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_23_321 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_35_192 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_50_151 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_11_505 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_23_365 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_1422_ _1422_/A1 _1569_/A2 _1569_/B1 _2171_/Q hold187/X vssd1 vssd1 vccd1 vccd1 _1422_/X
+ sky130_fd_sc_hd__a221o_1
XANTENNA__1326__B2 _2203_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_1353_ input16/X _1533_/A2 _1529_/B1 _2194_/Q hold244/X vssd1 vssd1 vccd1 vccd1 _1353_/X
+ sky130_fd_sc_hd__a221o_1
XANTENNA__1903__A _1913_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_1284_ input41/X _1529_/A2 _1529_/B1 _2217_/Q hold401/X vssd1 vssd1 vccd1 vccd1 _1284_/X
+ sky130_fd_sc_hd__a221o_1
XANTENNA__1629__A2 _1637_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_58_251 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_46_468 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_33_107 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_33_118 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_0999_ hold21/X _1012_/D _1012_/C _1012_/B vssd1 vssd1 vccd1 vccd1 hold22/A sky130_fd_sc_hd__and4b_1
XFILLER_0_26_170 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_41_140 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__1565__B2 _2104_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_14_376 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_1_281 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__1317__B2 _2206_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_9_381 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_24_107 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__1707__B _1761_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__1308__B2 _2209_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_46_38 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XANTENNA__1723__A _2151_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_1971_ _1979_/A vssd1 vssd1 vccd1 vccd1 _1971_/Y sky130_fd_sc_hd__inv_2
XFILLER_0_43_449 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__1547__B2 _2113_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__1547__A1 _1547_/A1 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_23_195 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_1405_ hold86/X hold949/X _1435_/S vssd1 vssd1 vccd1 vccd1 _2176_/D sky130_fd_sc_hd__mux2_1
X_1336_ hold337/X hold968/X hold27/X vssd1 vssd1 vccd1 vccd1 _2199_/D sky130_fd_sc_hd__mux2_1
Xinput1 data_in[0] vssd1 vssd1 vccd1 vccd1 input1/X sky130_fd_sc_hd__buf_1
X_1267_ hold501/X _2222_/Q hold26/X vssd1 vssd1 vccd1 vccd1 _1267_/X sky130_fd_sc_hd__mux2_1
X_1198_ _1198_/A _1198_/B _1198_/C vssd1 vssd1 vccd1 vccd1 _1198_/X sky130_fd_sc_hd__and3_1
XANTENNA__1483__B1 _1503_/B1 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_19_413 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_46_265 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_34_405 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_34_416 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_15_641 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__1538__A1 _2117_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_30_633 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
Xoutput360 _1682_/X vssd1 vssd1 vccd1 vccd1 data_out[40] sky130_fd_sc_hd__buf_12
Xoutput371 _1692_/X vssd1 vssd1 vccd1 vccd1 data_out[50] sky130_fd_sc_hd__buf_12
XFILLER_0_30_699 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xoutput382 _1702_/X vssd1 vssd1 vccd1 vccd1 data_out[60] sky130_fd_sc_hd__buf_12
Xoutput393 _1712_/X vssd1 vssd1 vccd1 vccd1 data_out[70] sky130_fd_sc_hd__buf_12
XFILLER_0_16_19 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_37_254 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_52_246 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__1529__A1 _1529_/A1 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_817 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_806 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_839 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_828 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_2170_ _2177_/CLK _2170_/D _1910_/Y vssd1 vssd1 vccd1 vccd1 _2170_/Q sky130_fd_sc_hd__dfrtp_4
X_1121_ hold643/X _1189_/A2 _1189_/B1 _1120_/X vssd1 vssd1 vccd1 vccd1 _2284_/D sky130_fd_sc_hd__a22o_1
X_1052_ _2230_/Q _2138_/Q _1094_/S vssd1 vssd1 vccd1 vccd1 _1052_/X sky130_fd_sc_hd__mux2_1
XFILLER_0_29_711 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_56_530 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_1954_ _1954_/A vssd1 vssd1 vccd1 vccd1 _1954_/Y sky130_fd_sc_hd__inv_2
XFILLER_0_16_416 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_28_243 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_28_265 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_43_213 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_1885_ _2039_/A vssd1 vssd1 vccd1 vccd1 _1885_/Y sky130_fd_sc_hd__inv_2
XFILLER_0_43_268 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_43_257 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_3_343 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_3_332 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_24_471 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_11_143 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_44_3 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_1319_ _1349_/A hold71/X vssd1 vssd1 vccd1 vccd1 hold72/A sky130_fd_sc_hd__and2_1
X_2299_ _2315_/CLK _2299_/D _2038_/Y vssd1 vssd1 vccd1 vccd1 _2299_/Q sky130_fd_sc_hd__dfrtp_1
XPHY_116 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_105 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_35_703 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_42_290 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__1392__C1 _1391_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XPHY_7 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_38_530 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_38_574 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_25_213 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_4_107 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_25_246 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_1670_ _2098_/Q _1677_/B vssd1 vssd1 vccd1 vccd1 _1670_/X sky130_fd_sc_hd__and2_1
XFILLER_0_40_227 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
Xhold309 _1508_/X vssd1 vssd1 vccd1 vccd1 _2132_/D sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA__1383__C1 hold529/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_603 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_614 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_625 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_658 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_636 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_647 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_2222_ _2225_/CLK _2222_/D _1962_/Y vssd1 vssd1 vccd1 vccd1 _2222_/Q sky130_fd_sc_hd__dfrtp_2
XTAP_669 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_2153_ _2328_/CLK _2153_/D _1896_/Y vssd1 vssd1 vccd1 vccd1 _2153_/Q sky130_fd_sc_hd__dfrtp_1
X_1104_ _2204_/Q _2112_/Q _1188_/S vssd1 vssd1 vccd1 vccd1 _1104_/X sky130_fd_sc_hd__mux2_1
XANTENNA__1911__A _1913_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_16_7 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_2084_ _2106_/CLK _2084_/D _1827_/Y vssd1 vssd1 vccd1 vccd1 _2084_/Q sky130_fd_sc_hd__dfrtp_4
X_1035_ hold599/X _1057_/A2 _1095_/B1 _1034_/X vssd1 vssd1 vccd1 vccd1 _2327_/D sky130_fd_sc_hd__a22o_1
XFILLER_0_29_541 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_44_500 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_33_83 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_44_533 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_1937_ _1957_/A vssd1 vssd1 vccd1 vccd1 _1937_/Y sky130_fd_sc_hd__inv_2
XANTENNA__1358__A _1415_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_1868_ _1954_/A vssd1 vssd1 vccd1 vccd1 _1868_/Y sky130_fd_sc_hd__inv_2
XFILLER_0_16_268 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xinput81 data_in[25] vssd1 vssd1 vccd1 vccd1 input81/X sky130_fd_sc_hd__buf_1
Xinput70 data_in[162] vssd1 vssd1 vccd1 vccd1 input70/X sky130_fd_sc_hd__buf_1
Xhold810 _2314_/Q vssd1 vssd1 vccd1 vccd1 hold810/X sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_31_249 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
Xhold821 _2287_/Q vssd1 vssd1 vccd1 vccd1 hold821/X sky130_fd_sc_hd__dlygate4sd3_1
Xinput92 data_in[35] vssd1 vssd1 vccd1 vccd1 input92/X sky130_fd_sc_hd__buf_1
X_1799_ _2237_/Q _1802_/B vssd1 vssd1 vccd1 vccd1 _1799_/X sky130_fd_sc_hd__and2_1
Xhold832 _2267_/Q vssd1 vssd1 vccd1 vccd1 hold832/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold854 _2305_/Q vssd1 vssd1 vccd1 vccd1 hold854/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold843 _1411_/X vssd1 vssd1 vccd1 vccd1 _2174_/D sky130_fd_sc_hd__dlygate4sd3_1
Xhold898 la_data_in[3] vssd1 vssd1 vccd1 vccd1 hold898/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold887 la_data_in[37] vssd1 vssd1 vccd1 vccd1 hold887/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold865 _2279_/Q vssd1 vssd1 vccd1 vccd1 hold865/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold876 _2292_/Q vssd1 vssd1 vccd1 vccd1 hold876/X sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA__1374__C1 hold127/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_58_91 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA_fanout584_A _1201_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__1141__A2 _1189_/A2 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xclkbuf_leaf_8_wb_clk_i clkbuf_leaf_9_wb_clk_i/A vssd1 vssd1 vccd1 vccd1 _2219_/CLK
+ sky130_fd_sc_hd__clkbuf_16
XANTENNA__1032__S _1094_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_39_349 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_47_393 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_35_511 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__1601__B1 _1623_/B1 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_35_599 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_50_536 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_22_238 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XANTENNA_hold963_A _2088_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__1365__C1 hold237/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__1715__B _1715_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__1207__S _1252_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__1380__A2 _1529_/A2 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__1731__A _2169_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_45_308 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_38_360 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_5_405 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_53_374 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_41_525 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_5_449 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_1722_ _2150_/Q _1804_/B vssd1 vssd1 vccd1 vccd1 _1722_/X sky130_fd_sc_hd__and2_1
XFILLER_0_13_238 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xhold106 _1346_/X vssd1 vssd1 vccd1 vccd1 hold106/X sky130_fd_sc_hd__dlymetal6s2s_1
Xhold117 _1424_/X vssd1 vssd1 vccd1 vccd1 hold117/X sky130_fd_sc_hd__dlymetal6s2s_1
X_1653_ _2081_/Q _1725_/B vssd1 vssd1 vccd1 vccd1 _1653_/X sky130_fd_sc_hd__and2_1
Xhold139 hold151/X vssd1 vssd1 vccd1 vccd1 hold139/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold128 _1374_/X vssd1 vssd1 vccd1 vccd1 hold128/X sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA__1356__C1 hold276/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_21_260 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_400 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_1584_ _1583_/X hold927/X _1622_/S vssd1 vssd1 vccd1 vccd1 _1584_/X sky130_fd_sc_hd__mux2_1
Xfanout608 _2034_/A vssd1 vssd1 vccd1 vccd1 _2033_/A sky130_fd_sc_hd__buf_8
XTAP_411 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_422 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_433 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_444 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_455 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_466 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_2205_ _2269_/CLK hold46/X _1945_/Y vssd1 vssd1 vccd1 vccd1 _2205_/Q sky130_fd_sc_hd__dfrtp_4
XTAP_477 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_488 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_499 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__1123__A2 _1183_/A2 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_2136_ _2315_/CLK _2136_/D _1879_/Y vssd1 vssd1 vccd1 vccd1 _2136_/Q sky130_fd_sc_hd__dfrtp_1
XFILLER_0_44_71 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_2067_ _2069_/A vssd1 vssd1 vccd1 vccd1 _2067_/Y sky130_fd_sc_hd__inv_2
X_1018_ _0972_/X hold36/X _0973_/B _0971_/C vssd1 vssd1 vccd1 vccd1 _1018_/Y sky130_fd_sc_hd__a211oi_1
XFILLER_0_29_382 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_29_393 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__1595__C1 _1391_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__1347__C1 hold106/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xhold662 hold805/X vssd1 vssd1 vccd1 vccd1 hold662/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold651 hold663/X vssd1 vssd1 vccd1 vccd1 hold651/X sky130_fd_sc_hd__dlymetal6s2s_1
Xhold640 hold693/X vssd1 vssd1 vccd1 vccd1 hold640/X sky130_fd_sc_hd__clkbuf_2
XFILLER_0_40_580 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xhold695 hold907/X vssd1 vssd1 vccd1 vccd1 hold695/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold684 hold810/X vssd1 vssd1 vccd1 vccd1 hold684/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold673 hold795/X vssd1 vssd1 vccd1 vccd1 hold673/X sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA__1362__A2 _1529_/A2 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_24_19 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_39_113 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_23_503 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_23_536 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_23_547 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__1726__A _2164_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_10_219 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xinput260 next_key vssd1 vssd1 vccd1 vccd1 _1202_/A2 sky130_fd_sc_hd__clkbuf_2
XFILLER_0_45_127 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_14_85 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_26_341 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_54_661 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_1705_ _2133_/Q _1724_/B vssd1 vssd1 vccd1 vccd1 _1705_/X sky130_fd_sc_hd__and2_1
XANTENNA__1577__C1 hold237/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_41_399 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_1636_ _1807_/A _1636_/B vssd1 vssd1 vccd1 vccd1 _2161_/D sky130_fd_sc_hd__nor2_1
X_1567_ input89/X _1569_/A2 _1569_/B1 _2103_/Q hold406/X vssd1 vssd1 vccd1 vccd1 _1567_/X
+ sky130_fd_sc_hd__a221o_1
XTAP_241 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_230 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_274 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_263 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_252 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_1498_ hold380/X _2137_/Q _1504_/S vssd1 vssd1 vccd1 vccd1 _1498_/X sky130_fd_sc_hd__mux2_1
XTAP_285 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_296 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_clkbuf_leaf_0_wb_clk_i_A clkbuf_leaf_9_wb_clk_i/A vssd1 vssd1 vccd1 vccd1
+ sky130_fd_sc_hd__diode_2
X_2119_ _2212_/CLK _2119_/D _1862_/Y vssd1 vssd1 vccd1 vccd1 _2119_/Q sky130_fd_sc_hd__dfrtp_4
XANTENNA_fanout547_A _1761_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_49_422 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_49_466 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_37_617 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_17_363 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_32_300 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_20_506 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_20_528 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_20_539 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_32_377 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__1583__A2 _1623_/A2 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xhold481 _1480_/X vssd1 vssd1 vccd1 vccd1 _2146_/D sky130_fd_sc_hd__dlygate4sd3_1
Xhold470 _1271_/X vssd1 vssd1 vccd1 vccd1 hold470/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold492 _0967_/Y vssd1 vssd1 vccd1 vccd1 _0973_/D sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA_hold926_A _2189_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_27_116 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_36_661 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_50_141 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_50_130 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_2_216 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_1421_ _1445_/A _1421_/B vssd1 vssd1 vccd1 vccd1 _1421_/X sky130_fd_sc_hd__and2_1
XANTENNA__1326__A2 _1197_/D vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_1352_ _1415_/A _1352_/B vssd1 vssd1 vccd1 vccd1 _1352_/X sky130_fd_sc_hd__and2_1
XANTENNA__1191__A hold38/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_1283_ _1310_/A _1283_/B vssd1 vssd1 vccd1 vccd1 _1283_/X sky130_fd_sc_hd__and2_1
XFILLER_0_25_84 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_18_138 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_42_631 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_0998_ _1014_/C _0997_/X _0995_/X _1197_/C vssd1 vssd1 vccd1 vccd1 _1192_/B sky130_fd_sc_hd__a211oi_4
Xclkbuf_leaf_22_wb_clk_i clkbuf_1_1__f_wb_clk_i/X vssd1 vssd1 vccd1 vccd1 _2291_/CLK
+ sky130_fd_sc_hd__clkbuf_16
XANTENNA__1565__A2 _1569_/A2 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xoutput520 _2247_/Q vssd1 vssd1 vccd1 vccd1 trigLoad sky130_fd_sc_hd__buf_12
X_1619_ _1619_/A1 _1619_/A2 _1619_/B1 _2077_/Q hold64/X vssd1 vssd1 vccd1 vccd1 _1619_/X
+ sky130_fd_sc_hd__a221o_1
XANTENNA__1317__A2 _1527_/A2 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__1040__S _1094_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_49_296 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_52_417 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_45_491 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__1308__A2 _1197_/D vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_1970_ _1979_/A vssd1 vssd1 vccd1 vccd1 _1970_/Y sky130_fd_sc_hd__inv_2
XFILLER_0_28_458 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_11_20 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_3_558 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__1547__A2 _1637_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_1404_ _1404_/A1 _1569_/A2 _1569_/B1 _2177_/Q hold85/X vssd1 vssd1 vccd1 vccd1 hold86/A
+ sky130_fd_sc_hd__a221o_1
XANTENNA__1180__A0 hold979/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_1335_ input22/X _1533_/A2 _1533_/B1 _2200_/Q hold336/X vssd1 vssd1 vccd1 vccd1 _1335_/X
+ sky130_fd_sc_hd__a221o_1
Xinput2 data_in[100] vssd1 vssd1 vccd1 vccd1 input2/X sky130_fd_sc_hd__clkbuf_1
X_1266_ input48/X _1519_/A2 _1519_/B1 _2223_/Q hold500/X vssd1 vssd1 vccd1 vccd1 _1266_/X
+ sky130_fd_sc_hd__a221o_1
X_1197_ _1197_/A _1197_/B _1197_/C _1197_/D vssd1 vssd1 vccd1 vccd1 _1197_/X sky130_fd_sc_hd__or4_1
XFILLER_0_36_83 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__1483__A1 _1483_/A1 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_59_561 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_52_60 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_46_211 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_19_447 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_15_620 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_14_163 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_30_645 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
Xoutput361 _1683_/X vssd1 vssd1 vccd1 vccd1 data_out[41] sky130_fd_sc_hd__buf_12
Xoutput350 _1673_/X vssd1 vssd1 vccd1 vccd1 data_out[31] sky130_fd_sc_hd__buf_12
XFILLER_0_30_678 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xoutput383 _1703_/X vssd1 vssd1 vccd1 vccd1 data_out[61] sky130_fd_sc_hd__buf_12
Xoutput394 _1713_/X vssd1 vssd1 vccd1 vccd1 data_out[71] sky130_fd_sc_hd__buf_12
Xoutput372 _1693_/X vssd1 vssd1 vccd1 vccd1 data_out[51] sky130_fd_sc_hd__buf_12
XANTENNA__1171__B1 _1189_/B1 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_37_222 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_18_480 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_25_417 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XANTENNA_hold993_A _2078_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__1718__B _1761_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_21_612 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__1529__A2 _1529_/A2 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_807 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__1734__A _2172_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_829 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_818 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_20_177 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_20_188 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_1120_ _2196_/Q _2104_/Q _1178_/S vssd1 vssd1 vccd1 vccd1 _1120_/X sky130_fd_sc_hd__mux2_1
XANTENNA__1162__A0 _2175_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_1051_ hold592/X _1057_/A2 _1057_/B1 _1050_/X vssd1 vssd1 vccd1 vccd1 _2319_/D sky130_fd_sc_hd__a22o_1
XFILLER_0_28_211 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_22_52 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_1953_ _1954_/A vssd1 vssd1 vccd1 vccd1 _1953_/Y sky130_fd_sc_hd__inv_2
XFILLER_0_56_586 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__1909__A _1922_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_1884_ _2039_/A vssd1 vssd1 vccd1 vccd1 _1884_/Y sky130_fd_sc_hd__inv_2
XFILLER_0_43_225 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_16_428 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_22_85 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_28_277 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_3_322 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_3_355 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_24_483 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_24_494 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__1644__A _2072_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_47_71 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__1153__B1 _1157_/B1 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_37_3 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_1318_ hold45/X _2205_/Q _1318_/S vssd1 vssd1 vccd1 vccd1 hold46/A sky130_fd_sc_hd__mux2_1
X_2298_ _2315_/CLK _2298_/D _2037_/Y vssd1 vssd1 vccd1 vccd1 _2298_/Q sky130_fd_sc_hd__dfrtp_1
X_1249_ hold313/X _2228_/Q _1252_/S vssd1 vssd1 vccd1 vccd1 _1249_/X sky130_fd_sc_hd__mux2_1
XANTENNA__1810__C _1810_/C vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_39_509 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XPHY_106 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_59_391 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XPHY_117 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_47_564 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_34_203 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_34_236 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_15_461 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XANTENNA__1392__B1 _1569_/B1 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__1144__A0 _2184_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__1447__A1 _2162_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XPHY_8 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__1729__A _2167_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_21_464 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_0_369 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_21_486 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_604 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_615 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_2221_ _2225_/CLK _2221_/D _1961_/Y vssd1 vssd1 vccd1 vccd1 _2221_/Q sky130_fd_sc_hd__dfrtp_4
XTAP_659 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_648 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_637 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_626 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__1135__B1 _1183_/B1 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_2152_ _2328_/CLK _2152_/D _1895_/Y vssd1 vssd1 vccd1 vccd1 _2152_/Q sky130_fd_sc_hd__dfrtp_1
XFILLER_0_17_41 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_1103_ hold593/X _1139_/A2 _1139_/B1 _1102_/X vssd1 vssd1 vccd1 vccd1 _2293_/D sky130_fd_sc_hd__a22o_1
XFILLER_0_17_63 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_2083_ _2106_/CLK _2083_/D _1826_/Y vssd1 vssd1 vccd1 vccd1 _2083_/Q sky130_fd_sc_hd__dfrtp_4
XFILLER_0_17_85 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__1438__A1 _2165_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_1034_ _2239_/Q _2147_/Q _1094_/S vssd1 vssd1 vccd1 vccd1 _1034_/X sky130_fd_sc_hd__mux2_1
XFILLER_0_56_350 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_16_203 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_16_214 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_1936_ _1957_/A vssd1 vssd1 vccd1 vccd1 _1936_/Y sky130_fd_sc_hd__inv_2
X_1867_ _1954_/A vssd1 vssd1 vccd1 vccd1 _1867_/Y sky130_fd_sc_hd__inv_2
XFILLER_0_44_589 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_4_642 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__1610__A1 _2081_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xinput82 data_in[26] vssd1 vssd1 vccd1 vccd1 input82/X sky130_fd_sc_hd__clkbuf_1
Xinput71 data_in[16] vssd1 vssd1 vccd1 vccd1 input71/X sky130_fd_sc_hd__clkbuf_1
Xinput60 data_in[153] vssd1 vssd1 vccd1 vccd1 input60/X sky130_fd_sc_hd__buf_1
X_1798_ _2236_/Q _1798_/B vssd1 vssd1 vccd1 vccd1 _1798_/X sky130_fd_sc_hd__and2_1
Xhold800 _2266_/Q vssd1 vssd1 vccd1 vccd1 hold800/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold811 _2256_/Q vssd1 vssd1 vccd1 vccd1 hold811/X sky130_fd_sc_hd__dlygate4sd3_1
Xinput93 data_in[36] vssd1 vssd1 vccd1 vccd1 input93/X sky130_fd_sc_hd__clkbuf_1
Xhold833 _2318_/Q vssd1 vssd1 vccd1 vccd1 hold833/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold844 la_data_in[43] vssd1 vssd1 vccd1 vccd1 hold844/X sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_12_442 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
Xhold855 _2278_/Q vssd1 vssd1 vccd1 vccd1 hold855/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold822 _2286_/Q vssd1 vssd1 vccd1 vccd1 hold822/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold866 _2329_/Q vssd1 vssd1 vccd1 vccd1 hold866/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold877 _2277_/Q vssd1 vssd1 vccd1 vccd1 hold877/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold888 _1558_/X vssd1 vssd1 vccd1 vccd1 _2107_/D sky130_fd_sc_hd__dlygate4sd3_1
Xhold899 _1438_/X vssd1 vssd1 vccd1 vccd1 _2165_/D sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA__1126__A0 _2193_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout577_A _1527_/B1 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__1429__A1 _2168_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_47_361 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_35_501 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__1601__B2 _2086_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_hold956_A _2097_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_38_29 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__1117__B1 _1183_/B1 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_26_512 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_5_417 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_26_556 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_38_394 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_1721_ _2149_/Q _1804_/B vssd1 vssd1 vccd1 vccd1 _1721_/X sky130_fd_sc_hd__and2_2
XFILLER_0_26_589 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_53_386 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
Xhold107 _1347_/X vssd1 vssd1 vccd1 vccd1 hold107/X sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_41_537 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_1652_ _2080_/Q _1725_/B vssd1 vssd1 vccd1 vccd1 _1652_/X sky130_fd_sc_hd__and2_1
Xhold118 _1425_/X vssd1 vssd1 vccd1 vccd1 hold118/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold129 _1375_/X vssd1 vssd1 vccd1 vccd1 _2186_/D sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA__1356__B1 _1529_/B1 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_1583_ input80/X _1623_/A2 _1623_/B1 _2095_/Q hold127/X vssd1 vssd1 vccd1 vccd1 _1583_/X
+ sky130_fd_sc_hd__a221o_1
Xfanout609 _2026_/A vssd1 vssd1 vccd1 vccd1 _2034_/A sky130_fd_sc_hd__clkbuf_8
XFILLER_0_21_294 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_401 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_412 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_423 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_434 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_445 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__1108__A0 _2202_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_456 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_467 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__1922__A _1922_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_2204_ _2269_/CLK hold74/X _1944_/Y vssd1 vssd1 vccd1 vccd1 _2204_/Q sky130_fd_sc_hd__dfrtp_4
XTAP_478 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_28_51 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_489 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__1641__B _1810_/C vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_2135_ _2239_/CLK _2135_/D _1878_/Y vssd1 vssd1 vccd1 vccd1 _2135_/Q sky130_fd_sc_hd__dfrtp_1
X_2066_ _2069_/A vssd1 vssd1 vccd1 vccd1 _2066_/Y sky130_fd_sc_hd__inv_2
X_1017_ _0983_/Y _1014_/C _0973_/B vssd1 vssd1 vccd1 vccd1 _1017_/X sky130_fd_sc_hd__o21ba_1
XFILLER_0_36_309 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_57_670 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_17_501 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_17_523 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_1919_ _1941_/A vssd1 vssd1 vccd1 vccd1 _1919_/Y sky130_fd_sc_hd__inv_2
XFILLER_0_17_567 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__1595__B1 _1623_/B1 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_8_61 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
Xhold630 hold737/X vssd1 vssd1 vccd1 vccd1 hold630/X sky130_fd_sc_hd__buf_1
XFILLER_0_12_250 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
Xhold663 hold848/X vssd1 vssd1 vccd1 vccd1 hold663/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold652 hold673/X vssd1 vssd1 vccd1 vccd1 hold652/X sky130_fd_sc_hd__clkbuf_2
Xhold641 hold682/X vssd1 vssd1 vccd1 vccd1 hold641/X sky130_fd_sc_hd__clkbuf_2
Xhold696 hold829/X vssd1 vssd1 vccd1 vccd1 hold696/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold674 hold853/X vssd1 vssd1 vccd1 vccd1 hold674/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold685 hold849/X vssd1 vssd1 vccd1 vccd1 hold685/X sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA__1832__A _1922_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_39_169 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_50_334 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__1742__A _2180_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xinput250 hold545/X vssd1 vssd1 vccd1 vccd1 _1453_/C sky130_fd_sc_hd__buf_1
Xinput261 slv_done vssd1 vssd1 vccd1 vccd1 _1637_/A sky130_fd_sc_hd__buf_2
XFILLER_0_14_20 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_45_106 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_18_309 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_45_139 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_5_225 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_26_353 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_1704_ _2132_/Q _1715_/B vssd1 vssd1 vccd1 vccd1 _1704_/X sky130_fd_sc_hd__and2_1
XFILLER_0_53_161 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_26_386 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_30_74 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__1917__A _1941_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_53_194 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_30_85 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_1635_ _1809_/B _1635_/B _1635_/C _1635_/D vssd1 vssd1 vccd1 vccd1 _1636_/B sky130_fd_sc_hd__or4_1
XANTENNA__1329__B1 _1541_/B1 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_1566_ _1565_/X hold933/X hold81/X vssd1 vssd1 vccd1 vccd1 _1566_/X sky130_fd_sc_hd__mux2_1
XFILLER_0_39_50 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_242 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_231 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_220 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_275 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_264 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_253 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__1652__A _2080_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_1497_ _1497_/A1 _1463_/B _1499_/B1 _2138_/Q hold379/X vssd1 vssd1 vccd1 vccd1 _1497_/X
+ sky130_fd_sc_hd__a221o_1
XTAP_286 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_297 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__1501__B1 _1503_/B1 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_2118_ _2212_/CLK _2118_/D _1861_/Y vssd1 vssd1 vccd1 vccd1 _2118_/Q sky130_fd_sc_hd__dfrtp_4
X_2049_ _2061_/A vssd1 vssd1 vccd1 vccd1 _2049_/Y sky130_fd_sc_hd__inv_2
XFILLER_0_36_128 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__1038__S _1038_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xhold460 _1484_/X vssd1 vssd1 vccd1 vccd1 _2144_/D sky130_fd_sc_hd__dlygate4sd3_1
Xhold471 _1515_/X vssd1 vssd1 vccd1 vccd1 hold471/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold493 _0973_/X vssd1 vssd1 vccd1 vccd1 hold493/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold482 la_data_in[58] vssd1 vssd1 vccd1 vccd1 hold482/X sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA__1099__A2 _1157_/A2 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_36_673 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__1559__B1 _1623_/B1 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_23_301 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__1737__A _2175_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_output361_A _1683_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_1420_ _1419_/X _2171_/Q hold27/X vssd1 vssd1 vccd1 vccd1 _1420_/X sky130_fd_sc_hd__mux2_1
X_1351_ _1350_/X hold959/X _1435_/S vssd1 vssd1 vccd1 vccd1 _1351_/X sky130_fd_sc_hd__mux2_1
X_1282_ _1281_/X _2217_/Q hold26/X vssd1 vssd1 vccd1 vccd1 _1282_/X sky130_fd_sc_hd__mux2_1
XFILLER_0_58_231 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_25_96 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__1411__S hold27/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_46_459 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_41_40 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_27_673 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__1647__A _2075_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_42_610 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_0997_ _0953_/Y _0992_/B _0990_/A _0991_/X _0959_/Y vssd1 vssd1 vccd1 vccd1 _0997_/X
+ sky130_fd_sc_hd__a32o_2
XFILLER_0_14_301 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_42_643 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xoutput510 hold578/X vssd1 vssd1 vccd1 vccd1 la_data_out[95] sky130_fd_sc_hd__buf_12
XFILLER_0_41_164 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_1618_ _1617_/X _2077_/Q _1622_/S vssd1 vssd1 vccd1 vccd1 _1618_/X sky130_fd_sc_hd__mux2_1
XFILLER_0_10_584 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_1549_ input99/X _1637_/B _1635_/C _2112_/Q hold183/X vssd1 vssd1 vccd1 vccd1 _1549_/X
+ sky130_fd_sc_hd__a221o_1
XFILLER_0_49_242 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__1321__S hold27/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_52_407 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_33_643 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_20_348 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_32_197 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_20_359 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__1292__A _1310_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xhold290 _1358_/X vssd1 vssd1 vccd1 vccd1 hold290/X sky130_fd_sc_hd__dlymetal6s2s_1
XANTENNA__1477__C1 hold298/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__1231__S _1252_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_55_223 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_28_426 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_43_429 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_3_537 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_24_643 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__1401__C1 hold132/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_24_687 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_11_348 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_1403_ _1415_/A hold84/X vssd1 vssd1 vccd1 vccd1 hold85/A sky130_fd_sc_hd__and2_1
XANTENNA__1633__C _1811_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_1334_ _1349_/A _1334_/B vssd1 vssd1 vccd1 vccd1 _1334_/X sky130_fd_sc_hd__and2_1
X_1265_ _1271_/A _1265_/B vssd1 vssd1 vccd1 vccd1 _1265_/X sky130_fd_sc_hd__and2_1
Xinput3 data_in[101] vssd1 vssd1 vccd1 vccd1 input3/X sky130_fd_sc_hd__clkbuf_1
XANTENNA__1930__A _1941_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_36_40 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_1196_ _2245_/Q _1200_/S hold549/X vssd1 vssd1 vccd1 vccd1 _1196_/X sky130_fd_sc_hd__a21o_1
XANTENNA__1483__A2 _1503_/A2 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_19_426 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_27_481 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_42_473 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_42_451 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_15_665 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_14_175 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_14_197 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_30_657 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xoutput340 _1664_/X vssd1 vssd1 vccd1 vccd1 data_out[22] sky130_fd_sc_hd__buf_12
Xoutput362 _1684_/X vssd1 vssd1 vccd1 vccd1 data_out[42] sky130_fd_sc_hd__buf_12
Xoutput351 _1674_/X vssd1 vssd1 vccd1 vccd1 data_out[32] sky130_fd_sc_hd__buf_12
XFILLER_0_2_592 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xoutput373 _1694_/X vssd1 vssd1 vccd1 vccd1 data_out[52] sky130_fd_sc_hd__buf_12
Xoutput395 _1714_/X vssd1 vssd1 vccd1 vccd1 data_out[72] sky130_fd_sc_hd__buf_12
Xoutput384 _1704_/X vssd1 vssd1 vccd1 vccd1 data_out[62] sky130_fd_sc_hd__buf_12
XANTENNA__1840__A _1922_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_37_234 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_37_278 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA_hold986_A _2185_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_33_462 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_808 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_819 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__1162__A1 _2083_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__1750__A _2188_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_clkbuf_leaf_24_wb_clk_i_A clkbuf_leaf_9_wb_clk_i/A vssd1 vssd1 vccd1 vccd1
+ sky130_fd_sc_hd__diode_2
X_1050_ _2231_/Q _2139_/Q _1094_/S vssd1 vssd1 vccd1 vccd1 _1050_/X sky130_fd_sc_hd__mux2_1
XANTENNA__1465__A2 _1466_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_1952_ _1954_/A vssd1 vssd1 vccd1 vccd1 _1952_/Y sky130_fd_sc_hd__inv_2
XFILLER_0_22_64 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_28_289 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_1883_ _1979_/A vssd1 vssd1 vccd1 vccd1 _1883_/Y sky130_fd_sc_hd__inv_2
XFILLER_0_24_462 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_51_281 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_3_367 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XANTENNA__1925__A _1941_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__1644__B _1725_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_47_61 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__1153__A1 hold570/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__1660__A _2088_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_2297_ _2330_/CLK _2297_/D _2036_/Y vssd1 vssd1 vccd1 vccd1 _2297_/Q sky130_fd_sc_hd__dfrtp_1
X_1317_ input29/X _1527_/A2 _1541_/B1 _2206_/Q hold44/X vssd1 vssd1 vccd1 vccd1 hold45/A
+ sky130_fd_sc_hd__a221o_1
X_1248_ input54/X _1463_/B _1499_/B1 _2229_/Q hold312/X vssd1 vssd1 vccd1 vccd1 _1248_/X
+ sky130_fd_sc_hd__a221o_1
XPHY_107 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_1179_ hold604/X _1189_/A2 _1189_/B1 _1178_/X vssd1 vssd1 vccd1 vccd1 _2255_/D sky130_fd_sc_hd__a22o_1
XPHY_118 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_19_201 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_47_554 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_19_234 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA_fanout522_A hold26/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_19_278 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_15_473 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__1835__A _1922_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_30_421 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_30_454 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__1392__B2 _2181_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__1046__S _1094_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__1144__A1 _2092_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XPHY_9 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__1729__B _1761_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_38_587 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_38_598 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XANTENNA__1080__A0 _2216_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_25_237 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__1745__A _2183_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_33_281 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_33_292 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__1383__B2 _2184_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_605 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_616 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_2220_ _2256_/CLK _2220_/D _1960_/Y vssd1 vssd1 vccd1 vccd1 _2220_/Q sky130_fd_sc_hd__dfrtp_4
XTAP_649 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_638 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_627 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_2151_ _2269_/CLK hold9/X _1894_/Y vssd1 vssd1 vccd1 vccd1 _2151_/Q sky130_fd_sc_hd__dfrtp_4
X_1102_ _2205_/Q _2113_/Q _1112_/S vssd1 vssd1 vccd1 vccd1 _1102_/X sky130_fd_sc_hd__mux2_1
X_2082_ _2106_/CLK _2082_/D _1825_/Y vssd1 vssd1 vccd1 vccd1 _2082_/Q sky130_fd_sc_hd__dfrtp_4
X_1033_ hold587/X _1057_/A2 _1057_/B1 _1032_/X vssd1 vssd1 vccd1 vccd1 _2328_/D sky130_fd_sc_hd__a22o_1
XFILLER_0_29_554 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_1935_ _1954_/A vssd1 vssd1 vccd1 vccd1 _1935_/Y sky130_fd_sc_hd__inv_2
XFILLER_0_8_459 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_44_546 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__1071__B1 _1097_/B1 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_1866_ _1954_/A vssd1 vssd1 vccd1 vccd1 _1866_/Y sky130_fd_sc_hd__inv_2
XFILLER_0_44_579 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_44_568 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
Xinput72 data_in[17] vssd1 vssd1 vccd1 vccd1 input72/X sky130_fd_sc_hd__buf_1
Xinput50 data_in[144] vssd1 vssd1 vccd1 vccd1 input50/X sky130_fd_sc_hd__buf_1
Xinput61 data_in[154] vssd1 vssd1 vccd1 vccd1 input61/X sky130_fd_sc_hd__dlymetal6s2s_1
X_1797_ _2235_/Q _1798_/B vssd1 vssd1 vccd1 vccd1 _1797_/X sky130_fd_sc_hd__and2_1
Xhold801 _2298_/Q vssd1 vssd1 vccd1 vccd1 hold801/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold812 _2299_/Q vssd1 vssd1 vccd1 vccd1 hold812/X sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA__1655__A _2083_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xinput94 data_in[37] vssd1 vssd1 vccd1 vccd1 input94/X sky130_fd_sc_hd__buf_1
Xinput83 data_in[27] vssd1 vssd1 vccd1 vccd1 input83/X sky130_fd_sc_hd__clkbuf_1
XFILLER_0_12_432 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
Xhold834 _2290_/Q vssd1 vssd1 vccd1 vccd1 hold834/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold845 _2317_/Q vssd1 vssd1 vccd1 vccd1 hold845/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold823 _2303_/Q vssd1 vssd1 vccd1 vccd1 hold823/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold867 _2250_/Q vssd1 vssd1 vccd1 vccd1 hold867/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold878 la_data_in[11] vssd1 vssd1 vccd1 vccd1 hold878/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold889 la_data_in[14] vssd1 vssd1 vccd1 vccd1 hold98/A sky130_fd_sc_hd__dlygate4sd3_1
Xhold856 _2281_/Q vssd1 vssd1 vccd1 vccd1 hold856/X sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA__1374__B2 _2187_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__1126__A1 _2101_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_47_384 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_35_535 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_35_557 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__1601__A2 _1623_/A2 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_22_207 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_15_281 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XANTENNA__1365__B2 _2190_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_hold949_A _2176_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__1504__S _1504_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_54_29 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_57_148 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_53_332 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_5_429 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_53_365 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_26_568 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_1720_ _2148_/Q _1802_/B vssd1 vssd1 vccd1 vccd1 _1720_/X sky130_fd_sc_hd__and2_1
XFILLER_0_53_398 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xhold108 la_data_in[94] vssd1 vssd1 vccd1 vccd1 hold108/X sky130_fd_sc_hd__dlygate4sd3_1
X_1651_ _2079_/Q _1725_/B vssd1 vssd1 vccd1 vccd1 _1651_/X sky130_fd_sc_hd__and2_1
Xhold119 hold507/X vssd1 vssd1 vccd1 vccd1 hold508/A sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA__1356__B2 _2193_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_1582_ hold209/X hold969/X _1622_/S vssd1 vssd1 vccd1 vccd1 _2095_/D sky130_fd_sc_hd__mux2_1
XTAP_402 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_413 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_424 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_435 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_446 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__1108__A1 _2110_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_457 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_2203_ _2251_/CLK _2203_/D _1943_/Y vssd1 vssd1 vccd1 vccd1 _2203_/Q sky130_fd_sc_hd__dfrtp_4
XTAP_479 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_468 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_28_74 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__1414__S hold27/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_28_85 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_2134_ _2239_/CLK _2134_/D _1877_/Y vssd1 vssd1 vccd1 vccd1 _2134_/Q sky130_fd_sc_hd__dfrtp_1
X_2065_ _2065_/A vssd1 vssd1 vccd1 vccd1 _2065_/Y sky130_fd_sc_hd__inv_2
X_1016_ hold110/X _1013_/X _0986_/A _0986_/B vssd1 vssd1 vccd1 vccd1 _1016_/X sky130_fd_sc_hd__a211o_1
Xclkbuf_leaf_16_wb_clk_i clkbuf_1_1__f_wb_clk_i/X vssd1 vssd1 vccd1 vccd1 _2296_/CLK
+ sky130_fd_sc_hd__clkbuf_16
XFILLER_0_9_713 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_8_234 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_8_223 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_29_373 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_44_365 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_1918_ _1941_/A vssd1 vssd1 vccd1 vccd1 _1918_/Y sky130_fd_sc_hd__inv_2
XFILLER_0_17_579 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__1595__B2 _2089_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_1849_ _1916_/A vssd1 vssd1 vccd1 vccd1 _1849_/Y sky130_fd_sc_hd__inv_2
Xhold620 hold661/X vssd1 vssd1 vccd1 vccd1 hold620/X sky130_fd_sc_hd__dlymetal6s2s_1
XANTENNA__1347__B2 _2196_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xhold653 hold715/X vssd1 vssd1 vccd1 vccd1 hold653/X sky130_fd_sc_hd__dlymetal6s2s_1
Xhold631 _1081_/X vssd1 vssd1 vccd1 vccd1 _2304_/D sky130_fd_sc_hd__dlygate4sd3_1
Xhold642 hold697/X vssd1 vssd1 vccd1 vccd1 hold642/X sky130_fd_sc_hd__clkbuf_2
Xhold675 hold851/X vssd1 vssd1 vccd1 vccd1 hold675/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold664 hold827/X vssd1 vssd1 vccd1 vccd1 hold664/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold697 hold820/X vssd1 vssd1 vccd1 vccd1 hold697/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold686 hold809/X vssd1 vssd1 vccd1 vccd1 hold686/X sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA__1324__S hold27/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_39_104 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_47_181 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_35_321 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__1035__B1 _1095_/B1 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_23_505 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_50_302 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_35_387 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__1295__A _1310_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__1338__B2 _2199_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__1234__S _1252_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xinput240 hold167/X vssd1 vssd1 vccd1 vccd1 hold168/A sky130_fd_sc_hd__clkbuf_1
Xinput251 hold426/X vssd1 vssd1 vccd1 vccd1 hold427/A sky130_fd_sc_hd__clkbuf_1
Xinput262 wb_rst_i vssd1 vssd1 vccd1 vccd1 input262/X sky130_fd_sc_hd__clkbuf_8
XFILLER_0_39_671 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_26_365 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_38_192 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_1703_ _2131_/Q _1715_/B vssd1 vssd1 vccd1 vccd1 _1703_/X sky130_fd_sc_hd__and2_1
XANTENNA__1577__B2 _2098_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_14_516 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_26_376 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_1634_ _1808_/C _1808_/D vssd1 vssd1 vccd1 vccd1 _1635_/D sky130_fd_sc_hd__nand2_1
XANTENNA__1329__B2 _2202_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_1565_ input90/X _1569_/A2 _1569_/B1 _2104_/Q hold106/X vssd1 vssd1 vccd1 vccd1 _1565_/X
+ sky130_fd_sc_hd__a221o_1
XTAP_232 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_210 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_221 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_265 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_254 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_243 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__1652__B _1725_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_1496_ _1495_/X _2138_/Q _1504_/S vssd1 vssd1 vccd1 vccd1 _1496_/X sky130_fd_sc_hd__mux2_1
XFILLER_0_39_95 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_287 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_276 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_298 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_55_50 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__1501__A1 _1501_/A1 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_55_83 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_2117_ _2173_/CLK _2117_/D _1860_/Y vssd1 vssd1 vccd1 vccd1 _2117_/Q sky130_fd_sc_hd__dfrtp_4
XFILLER_0_12_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_2048_ _2061_/A vssd1 vssd1 vccd1 vccd1 _2048_/Y sky130_fd_sc_hd__inv_2
XFILLER_0_49_457 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_17_310 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_17_343 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA_fanout602_A input262/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_44_195 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xhold472 _1516_/X vssd1 vssd1 vccd1 vccd1 _2128_/D sky130_fd_sc_hd__dlygate4sd3_1
Xhold461 hold466/X vssd1 vssd1 vccd1 vccd1 hold461/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold450 _1277_/X vssd1 vssd1 vccd1 vccd1 hold450/X sky130_fd_sc_hd__buf_1
Xhold483 _1273_/X vssd1 vssd1 vccd1 vccd1 _2220_/D sky130_fd_sc_hd__dlygate4sd3_1
Xhold494 _1020_/X vssd1 vssd1 vccd1 vccd1 hold494/X sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA__1054__S _1094_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__1559__B2 _2107_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_23_324 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_35_162 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_50_110 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_23_357 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_50_154 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_1350_ input17/X _1533_/A2 _1533_/B1 _2195_/Q hold406/X vssd1 vssd1 vccd1 vccd1 _1350_/X
+ sky130_fd_sc_hd__a221o_1
XANTENNA__1753__A _2191_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_1281_ input42/X _1527_/A2 _1527_/B1 _2218_/Q hold391/X vssd1 vssd1 vccd1 vccd1 _1281_/X
+ sky130_fd_sc_hd__a221o_1
XANTENNA__1928__A _1941_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_42_622 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_42_600 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_0996_ hold548/X hold759/X _0974_/X vssd1 vssd1 vccd1 vccd1 _0996_/X sky130_fd_sc_hd__o21a_1
XFILLER_0_14_313 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_54_493 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_42_699 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xoutput511 hold644/X vssd1 vssd1 vccd1 vccd1 la_data_out[96] sky130_fd_sc_hd__buf_12
Xoutput500 hold656/X vssd1 vssd1 vccd1 vccd1 la_data_out[85] sky130_fd_sc_hd__buf_12
XFILLER_0_14_379 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_1617_ _1617_/A1 _1619_/A2 _1619_/B1 _2078_/Q hold117/X vssd1 vssd1 vccd1 vccd1 _1617_/X
+ sky130_fd_sc_hd__a221o_1
XANTENNA__1663__A _2091_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_22_390 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_1548_ _1547_/X _2112_/Q _1632_/S vssd1 vssd1 vccd1 vccd1 _1548_/X sky130_fd_sc_hd__mux2_1
X_1479_ _1479_/A1 _1503_/A2 _1503_/B1 _2147_/Q hold415/X vssd1 vssd1 vccd1 vccd1 _1479_/X
+ sky130_fd_sc_hd__a221o_1
XANTENNA_fanout552_A _1157_/B1 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_37_416 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_9_351 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_9_340 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_37_449 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_18_663 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_45_482 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_45_471 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_32_154 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__1410__B1 _1201_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xhold280 hold280/A vssd1 vssd1 vccd1 vccd1 _1433_/B sky130_fd_sc_hd__dlygate4sd3_1
Xhold291 _1573_/X vssd1 vssd1 vccd1 vccd1 hold291/X sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA_hold931_A _2206_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_clkbuf_leaf_14_wb_clk_i_A clkbuf_1_1__f_wb_clk_i/X vssd1 vssd1 vccd1 vccd1
+ sky130_fd_sc_hd__diode_2
XANTENNA__1512__S _1520_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__1748__A _2186_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_23_110 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_23_132 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_23_165 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_24_677 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_24_699 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_1402_ hold133/X hold923/X _1435_/S vssd1 vssd1 vccd1 vccd1 _2177_/D sky130_fd_sc_hd__mux2_1
X_1333_ hold228/X hold948/X hold27/X vssd1 vssd1 vccd1 vccd1 _2200_/D sky130_fd_sc_hd__mux2_1
X_1264_ hold374/X hold924/X hold26/X vssd1 vssd1 vccd1 vccd1 _2223_/D sky130_fd_sc_hd__mux2_1
Xinput4 data_in[102] vssd1 vssd1 vccd1 vccd1 input4/X sky130_fd_sc_hd__clkbuf_1
XANTENNA__1468__B1 _1541_/B1 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_36_63 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_1195_ hold38/X _2246_/Q _1200_/S vssd1 vssd1 vccd1 vccd1 _1195_/X sky130_fd_sc_hd__mux2_1
XFILLER_0_59_530 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_19_449 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__1658__A _2086_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__1640__B1 _1637_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_6_365 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_0979_ _0979_/A _1453_/C vssd1 vssd1 vccd1 vccd1 _0980_/B sky130_fd_sc_hd__xor2_1
XFILLER_0_15_644 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_14_187 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xoutput352 _1675_/X vssd1 vssd1 vccd1 vccd1 data_out[33] sky130_fd_sc_hd__buf_12
Xoutput341 _1665_/X vssd1 vssd1 vccd1 vccd1 data_out[23] sky130_fd_sc_hd__buf_12
Xoutput330 _1802_/X vssd1 vssd1 vccd1 vccd1 data_out[160] sky130_fd_sc_hd__buf_12
Xoutput396 _1715_/X vssd1 vssd1 vccd1 vccd1 data_out[73] sky130_fd_sc_hd__buf_12
Xoutput363 _1685_/X vssd1 vssd1 vccd1 vccd1 data_out[43] sky130_fd_sc_hd__buf_12
Xoutput385 _1705_/X vssd1 vssd1 vccd1 vccd1 data_out[63] sky130_fd_sc_hd__buf_12
Xoutput374 _1695_/X vssd1 vssd1 vccd1 vccd1 data_out[53] sky130_fd_sc_hd__buf_12
XANTENNA__1171__A2 _1189_/A2 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__1459__B1 _1810_/C vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_25_408 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_52_249 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_33_430 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_33_474 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__1395__C1 _1394_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_hold979_A _2166_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_20_157 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_809 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__1750__B _1761_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xfanout590 _1038_/S vssd1 vssd1 vccd1 vccd1 _1094_/S sky130_fd_sc_hd__buf_6
XFILLER_0_29_703 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_28_246 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_1951_ _1954_/A vssd1 vssd1 vccd1 vccd1 _1951_/Y sky130_fd_sc_hd__inv_2
XFILLER_0_43_216 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_16_408 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_16_419 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_22_76 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_1882_ _1979_/A vssd1 vssd1 vccd1 vccd1 _1882_/Y sky130_fd_sc_hd__inv_2
XFILLER_0_24_441 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__1386__C1 hold521/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_51_260 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_3_379 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_51_293 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_11_135 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__1417__S hold27/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_1316_ _1349_/A hold43/X vssd1 vssd1 vccd1 vccd1 hold44/A sky130_fd_sc_hd__and2_1
XANTENNA__1941__A _1941_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__1153__A2 _1157_/A2 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_2296_ _2296_/CLK _2296_/D _2035_/Y vssd1 vssd1 vccd1 vccd1 _2296_/Q sky130_fd_sc_hd__dfrtp_1
X_1247_ _1271_/A _1247_/B vssd1 vssd1 vccd1 vccd1 _1247_/X sky130_fd_sc_hd__and2_1
X_1178_ _2167_/Q _2075_/Q _1178_/S vssd1 vssd1 vccd1 vccd1 _1178_/X sky130_fd_sc_hd__mux2_1
XPHY_119 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_108 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_47_533 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_47_522 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_47_511 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_35_706 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA_20 _2223_/CLK vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_34_249 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_42_293 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XANTENNA__1327__S hold27/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__1392__A2 _1569_/A2 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_30_499 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_38_522 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__1298__A _1310_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_38_533 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_53_503 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_53_558 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__1368__C1 hold248/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__1237__S _1252_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_21_444 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_21_455 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_606 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_617 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_639 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_628 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__1761__A _2199_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__1135__A2 _1157_/A2 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_2150_ _2322_/CLK _2150_/D _1893_/Y vssd1 vssd1 vccd1 vccd1 _2150_/Q sky130_fd_sc_hd__dfrtp_1
X_1101_ _2294_/Q _1139_/A2 _1139_/B1 _1100_/X vssd1 vssd1 vccd1 vccd1 _1101_/X sky130_fd_sc_hd__a22o_1
X_2081_ _2164_/CLK _2081_/D _1824_/Y vssd1 vssd1 vccd1 vccd1 _2081_/Q sky130_fd_sc_hd__dfrtp_4
X_1032_ _2240_/Q _2148_/Q _1094_/S vssd1 vssd1 vccd1 vccd1 _1032_/X sky130_fd_sc_hd__mux2_1
XFILLER_0_29_511 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_8_405 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_29_544 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_33_86 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_1934_ _1954_/A vssd1 vssd1 vccd1 vccd1 _1934_/Y sky130_fd_sc_hd__inv_2
XFILLER_0_44_514 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_29_577 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_44_536 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_16_249 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xinput40 data_in[135] vssd1 vssd1 vccd1 vccd1 input40/X sky130_fd_sc_hd__clkbuf_1
XANTENNA__1936__A _1957_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_32_709 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_1865_ _1954_/A vssd1 vssd1 vccd1 vccd1 _1865_/Y sky130_fd_sc_hd__inv_2
Xinput51 data_in[145] vssd1 vssd1 vccd1 vccd1 input51/X sky130_fd_sc_hd__buf_1
Xinput73 data_in[18] vssd1 vssd1 vccd1 vccd1 input73/X sky130_fd_sc_hd__clkbuf_1
Xinput62 data_in[155] vssd1 vssd1 vccd1 vccd1 input62/X sky130_fd_sc_hd__clkbuf_2
XANTENNA__1359__C1 hold290/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_1796_ _2234_/Q _1798_/B vssd1 vssd1 vccd1 vccd1 _1796_/X sky130_fd_sc_hd__and2_1
Xhold802 _2285_/Q vssd1 vssd1 vccd1 vccd1 hold802/X sky130_fd_sc_hd__dlygate4sd3_1
Xinput84 data_in[28] vssd1 vssd1 vccd1 vccd1 input84/X sky130_fd_sc_hd__clkbuf_1
Xinput95 data_in[38] vssd1 vssd1 vccd1 vccd1 input95/X sky130_fd_sc_hd__buf_1
Xhold835 _2252_/Q vssd1 vssd1 vccd1 vccd1 hold835/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold824 _2261_/Q vssd1 vssd1 vccd1 vccd1 hold824/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold846 _2295_/Q vssd1 vssd1 vccd1 vccd1 hold846/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold813 _2263_/Q vssd1 vssd1 vccd1 vccd1 hold813/X sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA__1655__B _1725_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xhold857 la_data_in[44] vssd1 vssd1 vccd1 vccd1 hold857/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold868 _2311_/Q vssd1 vssd1 vccd1 vccd1 hold868/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold879 _1414_/X vssd1 vssd1 vccd1 vccd1 _2173_/D sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_58_83 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__1671__A _2099_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_42_3 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_2279_ _2291_/CLK _2279_/D _2018_/Y vssd1 vssd1 vccd1 vccd1 _2279_/Q sky130_fd_sc_hd__dfrtp_1
XANTENNA__1610__S hold80/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__2007__A _2026_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_35_514 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_35_525 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_35_547 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_7_471 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_15_271 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_15_293 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__1365__A2 _1529_/A2 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__1117__A2 _1183_/A2 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__1520__S _1520_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__1589__C1 hold529/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__1756__A _2194_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_1650_ _2078_/Q _1677_/B vssd1 vssd1 vccd1 vccd1 _1650_/X sky130_fd_sc_hd__and2_1
XFILLER_0_34_580 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_1581_ input81/X _1623_/A2 _1623_/B1 _2096_/Q hold208/X vssd1 vssd1 vccd1 vccd1 _1581_/X
+ sky130_fd_sc_hd__a221o_1
Xhold109 hold109/A vssd1 vssd1 vccd1 vccd1 _1002_/A sky130_fd_sc_hd__clkbuf_2
XTAP_403 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_414 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_425 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_436 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_447 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_458 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_2202_ _2212_/CLK _2202_/D _1942_/Y vssd1 vssd1 vccd1 vccd1 _2202_/Q sky130_fd_sc_hd__dfrtp_4
XTAP_469 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_28_97 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_2133_ _2300_/CLK _2133_/D _1876_/Y vssd1 vssd1 vccd1 vccd1 _2133_/Q sky130_fd_sc_hd__dfrtp_1
XFILLER_0_44_52 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_2064_ _2069_/A vssd1 vssd1 vccd1 vccd1 _2064_/Y sky130_fd_sc_hd__inv_2
XFILLER_0_44_85 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_44_74 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_1015_ _1011_/X hold77/X _1192_/B vssd1 vssd1 vccd1 vccd1 hold78/A sky130_fd_sc_hd__o21a_1
XFILLER_0_29_330 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_44_322 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_29_385 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_29_396 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_1917_ _1941_/A vssd1 vssd1 vccd1 vccd1 _1917_/Y sky130_fd_sc_hd__inv_2
XANTENNA__1666__A _2094_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_44_377 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_1848_ _1916_/A vssd1 vssd1 vccd1 vccd1 _1848_/Y sky130_fd_sc_hd__inv_2
XFILLER_0_4_430 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_12_230 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xhold621 hold671/X vssd1 vssd1 vccd1 vccd1 hold621/X sky130_fd_sc_hd__buf_1
Xhold610 hold733/X vssd1 vssd1 vccd1 vccd1 hold610/X sky130_fd_sc_hd__buf_1
X_1779_ _2217_/Q _1798_/B vssd1 vssd1 vccd1 vccd1 _1779_/X sky130_fd_sc_hd__and2_1
Xhold654 _1087_/X vssd1 vssd1 vccd1 vccd1 _2301_/D sky130_fd_sc_hd__dlygate4sd3_1
Xhold643 hold662/X vssd1 vssd1 vccd1 vccd1 hold643/X sky130_fd_sc_hd__buf_1
Xhold632 hold695/X vssd1 vssd1 vccd1 vccd1 hold632/X sky130_fd_sc_hd__dlymetal6s2s_1
Xhold665 hold803/X vssd1 vssd1 vccd1 vccd1 hold665/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold676 hold852/X vssd1 vssd1 vccd1 vccd1 hold676/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold687 hold799/X vssd1 vssd1 vccd1 vccd1 hold687/X sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_40_583 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xhold698 hold847/X vssd1 vssd1 vccd1 vccd1 hold698/X sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_35_377 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_31_550 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_31_561 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XANTENNA_hold961_A _2201_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xinput230 hold62/X vssd1 vssd1 vccd1 vccd1 hold63/A sky130_fd_sc_hd__buf_1
Xinput241 hold115/X vssd1 vssd1 vccd1 vccd1 hold116/A sky130_fd_sc_hd__clkbuf_1
Xinput252 hold185/X vssd1 vssd1 vccd1 vccd1 hold186/A sky130_fd_sc_hd__buf_1
XFILLER_0_39_650 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_14_99 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_38_160 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_30_21 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_1702_ _2130_/Q _1715_/B vssd1 vssd1 vccd1 vccd1 _1702_/X sky130_fd_sc_hd__and2_1
XFILLER_0_30_43 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_1633_ hold2/A hold88/A _1811_/A _1025_/Y vssd1 vssd1 vccd1 vccd1 _1807_/A sky130_fd_sc_hd__or4b_2
XFILLER_0_10_701 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_1_411 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_1_444 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__1329__A2 _1197_/D vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_1564_ hold137/X hold940/X hold81/X vssd1 vssd1 vccd1 vccd1 _2104_/D sky130_fd_sc_hd__mux2_1
XTAP_233 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_211 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_222 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_200 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_1495_ _1495_/A1 _1495_/A2 _1495_/B1 _2139_/Q hold359/X vssd1 vssd1 vccd1 vccd1 _1495_/X
+ sky130_fd_sc_hd__a221o_1
XTAP_266 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_255 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_244 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_288 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_277 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_299 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__1501__A2 _1503_/A2 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_2116_ _2173_/CLK _2116_/D _1859_/Y vssd1 vssd1 vccd1 vccd1 _2116_/Q sky130_fd_sc_hd__dfrtp_4
XFILLER_0_49_425 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_49_414 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_2047_ _2065_/A vssd1 vssd1 vccd1 vccd1 _2047_/Y sky130_fd_sc_hd__inv_2
XFILLER_0_49_447 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_49_469 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_37_609 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_45_631 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_45_620 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_44_141 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_17_355 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xhold451 _1278_/X vssd1 vssd1 vccd1 vccd1 hold451/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold440 _1285_/X vssd1 vssd1 vccd1 vccd1 _2216_/D sky130_fd_sc_hd__dlygate4sd3_1
Xhold462 hold462/A vssd1 vssd1 vccd1 vccd1 _1268_/B sky130_fd_sc_hd__dlygate4sd3_1
Xhold495 _1190_/X vssd1 vssd1 vccd1 vccd1 _1191_/C sky130_fd_sc_hd__dlygate4sd3_1
Xhold473 hold478/X vssd1 vssd1 vccd1 vccd1 hold473/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold484 la_data_in[87] vssd1 vssd1 vccd1 vccd1 hold484/X sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_40_391 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_35_130 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__1559__A2 _1623_/A2 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_2_219 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_50_166 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_11_509 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xclkbuf_leaf_1_wb_clk_i clkbuf_leaf_9_wb_clk_i/A vssd1 vssd1 vccd1 vccd1 _2212_/CLK
+ sky130_fd_sc_hd__clkbuf_16
XFILLER_0_31_391 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_1280_ _1310_/A _1280_/B vssd1 vssd1 vccd1 vccd1 _1280_/X sky130_fd_sc_hd__and2_1
XANTENNA__1495__A1 _1495_/A1 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_25_43 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_58_211 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_46_439 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_27_620 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_6_536 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_39_491 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_0995_ _0978_/A _0978_/B _1012_/D _1012_/C vssd1 vssd1 vccd1 vccd1 _0995_/X sky130_fd_sc_hd__and4bb_2
XFILLER_0_26_141 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_41_86 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xoutput501 hold630/X vssd1 vssd1 vccd1 vccd1 la_data_out[86] sky130_fd_sc_hd__buf_12
XANTENNA__1944__A _1949_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xoutput512 hold573/X vssd1 vssd1 vccd1 vccd1 la_data_out[97] sky130_fd_sc_hd__buf_12
X_1616_ hold188/X hold993/X _1632_/S vssd1 vssd1 vccd1 vccd1 _2078_/D sky130_fd_sc_hd__mux2_1
XFILLER_0_10_531 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__1183__B1 _1183_/B1 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_1547_ _1547_/A1 _1637_/B _1635_/C _2113_/Q hold72/X vssd1 vssd1 vccd1 vccd1 _1547_/X
+ sky130_fd_sc_hd__a221o_1
X_1478_ hold299/X _2147_/Q _1504_/S vssd1 vssd1 vccd1 vccd1 _1478_/X sky130_fd_sc_hd__mux2_1
XFILLER_0_49_211 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_18_653 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_45_461 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_33_612 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_45_494 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__1410__B2 _2175_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_20_317 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
Xhold270 hold270/A vssd1 vssd1 vccd1 vccd1 _1205_/B sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA__1174__A0 _2169_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xhold292 la_data_in[52] vssd1 vssd1 vccd1 vccd1 hold292/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold281 _1433_/X vssd1 vssd1 vccd1 vccd1 hold281/X sky130_fd_sc_hd__buf_1
XANTENNA_hold924_A _2223_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__1477__A1 _1477_/A1 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_55_214 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__1748__B _1761_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_24_601 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_36_461 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_36_472 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_24_645 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XANTENNA__1401__B2 _2178_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__1764__A _2202_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_1401_ _1401_/A1 _1533_/A2 _1533_/B1 _2178_/Q hold132/X vssd1 vssd1 vccd1 vccd1 _1401_/X
+ sky130_fd_sc_hd__a221o_1
XANTENNA__1165__B1 _1183_/B1 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_1332_ input24/X _1197_/D _1541_/B1 _2201_/Q hold227/X vssd1 vssd1 vccd1 vccd1 _1332_/X
+ sky130_fd_sc_hd__a221o_1
X_1263_ input49/X _1519_/A2 _1519_/B1 _2224_/Q hold373/X vssd1 vssd1 vccd1 vccd1 _1263_/X
+ sky130_fd_sc_hd__a221o_1
Xinput5 data_in[103] vssd1 vssd1 vccd1 vccd1 input5/X sky130_fd_sc_hd__clkbuf_1
XANTENNA__1468__A1 _1310_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_1194_ _1194_/A _1194_/B _1193_/Y vssd1 vssd1 vccd1 vccd1 _1194_/X sky130_fd_sc_hd__or3b_1
XANTENNA__1468__B2 _2162_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_59_564 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_59_586 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_46_214 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_52_85 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_46_269 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_15_612 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_6_377 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_0978_ _0978_/A _0978_/B hold36/X vssd1 vssd1 vccd1 vccd1 _1453_/D sky130_fd_sc_hd__or3_1
XFILLER_0_15_623 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_15_656 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_15_689 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__1674__A _2102_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xoutput353 _1676_/X vssd1 vssd1 vccd1 vccd1 data_out[34] sky130_fd_sc_hd__buf_12
Xoutput342 _1666_/X vssd1 vssd1 vccd1 vccd1 data_out[24] sky130_fd_sc_hd__buf_12
Xoutput320 _1793_/X vssd1 vssd1 vccd1 vccd1 data_out[151] sky130_fd_sc_hd__buf_12
Xoutput331 _1803_/X vssd1 vssd1 vccd1 vccd1 data_out[161] sky130_fd_sc_hd__buf_12
Xoutput386 _1706_/X vssd1 vssd1 vccd1 vccd1 data_out[64] sky130_fd_sc_hd__buf_12
Xoutput364 _1686_/X vssd1 vssd1 vccd1 vccd1 data_out[44] sky130_fd_sc_hd__buf_12
Xoutput375 _1696_/X vssd1 vssd1 vccd1 vccd1 data_out[54] sky130_fd_sc_hd__buf_12
XANTENNA__1156__A0 _2178_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_10_372 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xoutput397 _1716_/X vssd1 vssd1 vccd1 vccd1 data_out[74] sky130_fd_sc_hd__buf_12
XFILLER_0_38_704 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_37_225 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__1631__A1 input1/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__1631__B2 _2071_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_33_442 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__1395__B1 _1569_/B1 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__1147__B1 _1189_/B1 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xfanout591 _1394_/A vssd1 vssd1 vccd1 vccd1 _1445_/A sky130_fd_sc_hd__buf_4
Xfanout580 _1201_/X vssd1 vssd1 vccd1 vccd1 _1527_/B1 sky130_fd_sc_hd__clkbuf_4
XANTENNA__1759__A _2197_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_28_214 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_7_119 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_1950_ _1954_/A vssd1 vssd1 vccd1 vccd1 _1950_/Y sky130_fd_sc_hd__inv_2
X_1881_ _1979_/A vssd1 vssd1 vccd1 vccd1 _1881_/Y sky130_fd_sc_hd__inv_2
XFILLER_0_36_291 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__1386__B1 _1529_/B1 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__1138__A0 _2187_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_1315_ hold198/X hold931/X _1318_/S vssd1 vssd1 vccd1 vccd1 _2206_/D sky130_fd_sc_hd__mux2_1
X_2295_ _2296_/CLK _2295_/D _2034_/Y vssd1 vssd1 vccd1 vccd1 _2295_/Q sky130_fd_sc_hd__dfrtp_1
X_1246_ _1245_/X _2229_/Q _1252_/S vssd1 vssd1 vccd1 vccd1 _1246_/X sky130_fd_sc_hd__mux2_1
X_1177_ hold658/X _1183_/A2 _1183_/B1 _1176_/X vssd1 vssd1 vccd1 vccd1 _2256_/D sky130_fd_sc_hd__a22o_1
XPHY_109 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__1669__A _2097_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_47_545 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_19_225 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_47_567 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_7_642 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA_10 la_data_in[53] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_21 hold42/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__1613__B2 _2080_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_42_272 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__1129__B1 _1189_/B1 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_38_501 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_38_545 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XANTENNA__1604__A1 _2084_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_hold991_A _2110_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__1518__S _1520_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_21_434 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_21_467 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_21_489 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_607 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_618 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_629 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__1761__B _1761_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_1100_ _2206_/Q _2114_/Q _1188_/S vssd1 vssd1 vccd1 vccd1 _1100_/X sky130_fd_sc_hd__mux2_1
XFILLER_0_17_55 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_2080_ _2164_/CLK hold56/X _1823_/Y vssd1 vssd1 vccd1 vccd1 _2080_/Q sky130_fd_sc_hd__dfrtp_4
X_1031_ hold588/X _1057_/A2 _1057_/B1 hold789/X vssd1 vssd1 vccd1 vccd1 _2329_/D sky130_fd_sc_hd__a22o_1
XFILLER_0_48_309 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_29_501 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_33_43 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_8_417 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_1933_ _1954_/A vssd1 vssd1 vccd1 vccd1 _1933_/Y sky130_fd_sc_hd__inv_2
XFILLER_0_33_98 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_16_217 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XANTENNA__1071__A2 _1097_/A2 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xinput30 data_in[126] vssd1 vssd1 vccd1 vccd1 input30/X sky130_fd_sc_hd__buf_1
XFILLER_0_44_559 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_1864_ _1954_/A vssd1 vssd1 vccd1 vccd1 _1864_/Y sky130_fd_sc_hd__inv_2
Xinput63 data_in[156] vssd1 vssd1 vccd1 vccd1 input63/X sky130_fd_sc_hd__clkbuf_2
Xinput52 data_in[146] vssd1 vssd1 vccd1 vccd1 input52/X sky130_fd_sc_hd__clkbuf_2
Xinput41 data_in[136] vssd1 vssd1 vccd1 vccd1 input41/X sky130_fd_sc_hd__clkbuf_1
XANTENNA__1359__B1 _1529_/B1 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_1795_ _2233_/Q _1798_/B vssd1 vssd1 vccd1 vccd1 _1795_/X sky130_fd_sc_hd__and2_1
Xhold803 _2330_/Q vssd1 vssd1 vccd1 vccd1 hold803/X sky130_fd_sc_hd__dlygate4sd3_1
Xinput85 data_in[29] vssd1 vssd1 vccd1 vccd1 input85/X sky130_fd_sc_hd__clkbuf_1
Xinput74 data_in[19] vssd1 vssd1 vccd1 vccd1 input74/X sky130_fd_sc_hd__clkbuf_1
Xinput96 data_in[39] vssd1 vssd1 vccd1 vccd1 input96/X sky130_fd_sc_hd__buf_1
Xhold836 _2273_/Q vssd1 vssd1 vccd1 vccd1 hold836/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold825 _2326_/Q vssd1 vssd1 vccd1 vccd1 hold825/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold814 _2296_/Q vssd1 vssd1 vccd1 vccd1 hold814/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold847 _2320_/Q vssd1 vssd1 vccd1 vccd1 hold847/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold869 la_data_in[40] vssd1 vssd1 vccd1 vccd1 hold869/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold858 _1544_/X vssd1 vssd1 vccd1 vccd1 _2114_/D sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_35_3 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_2278_ _2300_/CLK _2278_/D _2017_/Y vssd1 vssd1 vccd1 vccd1 _2278_/Q sky130_fd_sc_hd__dfrtp_1
X_1229_ _1277_/A _1229_/B vssd1 vssd1 vccd1 vccd1 _1229_/X sky130_fd_sc_hd__and2_1
XFILLER_0_47_397 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_50_529 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_43_592 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_30_242 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_30_253 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_30_286 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__1862__A _1941_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_38_320 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_53_312 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_26_515 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_38_375 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_1580_ _1579_/X hold938/X _1622_/S vssd1 vssd1 vccd1 vccd1 _1580_/X sky130_fd_sc_hd__mux2_1
XFILLER_0_21_297 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_404 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_415 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__1772__A _2210_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_426 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_437 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_448 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__1513__B1 _1519_/B1 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_459 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_2201_ _2212_/CLK _2201_/D _1941_/Y vssd1 vssd1 vccd1 vccd1 _2201_/Q sky130_fd_sc_hd__dfrtp_4
X_2132_ _2224_/CLK _2132_/D _1875_/Y vssd1 vssd1 vccd1 vccd1 _2132_/Q sky130_fd_sc_hd__dfrtp_1
X_2063_ _2069_/A vssd1 vssd1 vccd1 vccd1 _2063_/Y sky130_fd_sc_hd__inv_2
XFILLER_0_44_64 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_1014_ hold76/X _1014_/B _1014_/C _1014_/D vssd1 vssd1 vccd1 vccd1 hold77/A sky130_fd_sc_hd__nand4_1
XFILLER_0_48_139 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_57_673 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_56_172 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_44_312 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_17_526 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__1947__A _1949_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_44_334 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_1916_ _1916_/A vssd1 vssd1 vccd1 vccd1 _1916_/Y sky130_fd_sc_hd__inv_2
X_1847_ _1916_/A vssd1 vssd1 vccd1 vccd1 _1847_/Y sky130_fd_sc_hd__inv_2
XFILLER_0_32_518 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xhold600 hold741/X vssd1 vssd1 vccd1 vccd1 hold600/X sky130_fd_sc_hd__dlymetal6s2s_1
XFILLER_0_8_75 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xclkbuf_leaf_25_wb_clk_i clkbuf_leaf_9_wb_clk_i/A vssd1 vssd1 vccd1 vccd1 _2249_/CLK
+ sky130_fd_sc_hd__clkbuf_16
Xhold611 _1141_/X vssd1 vssd1 vccd1 vccd1 _2274_/D sky130_fd_sc_hd__dlygate4sd3_1
X_1778_ _2216_/Q _1798_/B vssd1 vssd1 vccd1 vccd1 _1778_/X sky130_fd_sc_hd__and2_1
XFILLER_0_12_253 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
Xhold633 hold734/X vssd1 vssd1 vccd1 vccd1 hold633/X sky130_fd_sc_hd__buf_1
Xhold622 _1109_/X vssd1 vssd1 vccd1 vccd1 _2290_/D sky130_fd_sc_hd__dlygate4sd3_1
Xhold644 hold684/X vssd1 vssd1 vccd1 vccd1 hold644/X sky130_fd_sc_hd__clkbuf_2
XFILLER_0_40_562 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__1682__A _2110_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xhold655 hold659/X vssd1 vssd1 vccd1 vccd1 hold655/X sky130_fd_sc_hd__clkbuf_2
Xhold677 hold846/X vssd1 vssd1 vccd1 vccd1 hold677/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold666 hold828/X vssd1 vssd1 vccd1 vccd1 hold666/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold688 hold796/X vssd1 vssd1 vccd1 vccd1 hold688/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold699 hold815/X vssd1 vssd1 vccd1 vccd1 hold699/X sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA_fanout575_A _1569_/B1 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__1857__A _1913_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_hold787_A _2211_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_31_573 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
Xinput220 hold498/X vssd1 vssd1 vccd1 vccd1 hold499/A sky130_fd_sc_hd__buf_1
Xinput231 hold408/X vssd1 vssd1 vccd1 vccd1 hold409/A sky130_fd_sc_hd__clkbuf_1
Xinput253 hold761/X vssd1 vssd1 vccd1 vccd1 _0992_/B sky130_fd_sc_hd__buf_1
Xinput242 hold269/X vssd1 vssd1 vccd1 vccd1 hold270/A sky130_fd_sc_hd__clkbuf_1
XFILLER_0_39_662 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__1767__A _2205_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_39_673 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_54_643 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_53_120 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_53_131 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_54_698 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_1701_ _2129_/Q _1715_/B vssd1 vssd1 vccd1 vccd1 _1701_/X sky130_fd_sc_hd__and2_1
XFILLER_0_41_304 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_53_197 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_41_337 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_1632_ hold50/X _2070_/Q _1632_/S vssd1 vssd1 vccd1 vccd1 hold51/A sky130_fd_sc_hd__mux2_1
X_1563_ input91/X _1569_/A2 _1569_/B1 _2105_/Q hold136/X vssd1 vssd1 vccd1 vccd1 _1563_/X
+ sky130_fd_sc_hd__a221o_1
XFILLER_0_10_713 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_212 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_223 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_201 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_1494_ hold437/X _2139_/Q _1504_/S vssd1 vssd1 vccd1 vccd1 _1494_/X sky130_fd_sc_hd__mux2_1
XFILLER_0_39_53 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_256 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_245 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_234 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_289 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_278 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_267 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__1441__S hold27/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_2115_ _2173_/CLK _2115_/D _1858_/Y vssd1 vssd1 vccd1 vccd1 _2115_/Q sky130_fd_sc_hd__dfrtp_4
X_2046_ _2065_/A vssd1 vssd1 vccd1 vccd1 _2046_/Y sky130_fd_sc_hd__inv_2
XANTENNA__1677__A _2105_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_29_172 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_17_334 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_29_183 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_17_378 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
Xhold430 _1016_/X vssd1 vssd1 vccd1 vccd1 hold430/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold452 la_data_in[56] vssd1 vssd1 vccd1 vccd1 hold452/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold441 hold459/X vssd1 vssd1 vccd1 vccd1 hold441/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold463 _1268_/X vssd1 vssd1 vccd1 vccd1 hold463/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold474 hold474/A vssd1 vssd1 vccd1 vccd1 _1256_/B sky130_fd_sc_hd__dlygate4sd3_1
Xhold485 _0979_/A vssd1 vssd1 vccd1 vccd1 _1453_/A sky130_fd_sc_hd__dlygate4sd3_1
Xhold496 hold780/X vssd1 vssd1 vccd1 vccd1 _2247_/D sky130_fd_sc_hd__dlygate4sd3_1
XTAP_790 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__1351__S _1435_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_48_470 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_36_698 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_50_134 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_23_337 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_50_145 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_50_178 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__1526__S hold80/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__1261__S hold26/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_59_713 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_58_278 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_41_54 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_42_613 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_0994_ hold783/X hold554/X _0974_/X hold37/X vssd1 vssd1 vccd1 vccd1 _0994_/X sky130_fd_sc_hd__o211a_1
XFILLER_0_26_197 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_41_101 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
Xoutput502 hold635/X vssd1 vssd1 vccd1 vccd1 la_data_out[87] sky130_fd_sc_hd__buf_12
XFILLER_0_41_167 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xoutput513 hold589/X vssd1 vssd1 vccd1 vccd1 la_data_out[98] sky130_fd_sc_hd__buf_12
XFILLER_0_1_220 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_1615_ _1615_/A1 _1623_/A2 _1635_/C _2079_/Q hold187/X vssd1 vssd1 vccd1 vccd1 _1615_/X
+ sky130_fd_sc_hd__a221o_1
X_1546_ _1545_/X hold797/X _1632_/S vssd1 vssd1 vccd1 vccd1 _2113_/D sky130_fd_sc_hd__mux2_1
XFILLER_0_10_587 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__1960__A _2002_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_1477_ _1477_/A1 _1495_/A2 _1495_/B1 _2148_/Q hold298/X vssd1 vssd1 vccd1 vccd1 _1477_/X
+ sky130_fd_sc_hd__a221o_1
X_2029_ _2033_/A vssd1 vssd1 vccd1 vccd1 _2029_/Y sky130_fd_sc_hd__inv_2
XANTENNA_fanout538_A _1520_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_49_289 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_18_643 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_17_142 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_17_164 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_18_687 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_17_197 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__1410__A2 _1569_/A2 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_20_329 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
Xhold271 _1205_/X vssd1 vssd1 vccd1 vccd1 hold271/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold260 la_data_in[31] vssd1 vssd1 vccd1 vccd1 hold260/X sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA__1174__A1 _2077_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xhold293 _1528_/X vssd1 vssd1 vccd1 vccd1 _2122_/D sky130_fd_sc_hd__dlygate4sd3_1
Xhold282 _1434_/X vssd1 vssd1 vccd1 vccd1 hold282/X sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA__1870__A _2002_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_28_418 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_28_429 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_24_613 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_36_451 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_23_123 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_24_657 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_24_668 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_23_189 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_1400_ _1415_/A _1400_/B vssd1 vssd1 vccd1 vccd1 _1400_/X sky130_fd_sc_hd__and2_1
X_1331_ _1349_/A _1331_/B vssd1 vssd1 vccd1 vccd1 _1331_/X sky130_fd_sc_hd__and2_1
XANTENNA__1780__A _2218_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_1262_ _1277_/A _1262_/B vssd1 vssd1 vccd1 vccd1 _1262_/X sky130_fd_sc_hd__and2_1
Xinput6 data_in[104] vssd1 vssd1 vccd1 vccd1 input6/X sky130_fd_sc_hd__clkbuf_1
X_1193_ _1810_/C _1805_/A vssd1 vssd1 vccd1 vccd1 _1193_/Y sky130_fd_sc_hd__nand2_4
XFILLER_0_52_97 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_6_312 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_54_281 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_54_270 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__1955__A _1957_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_0977_ hold35/X _0977_/B _0977_/C _0977_/D vssd1 vssd1 vccd1 vccd1 hold36/A sky130_fd_sc_hd__nand4_1
XFILLER_0_15_635 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_27_473 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_42_454 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_6_389 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_15_668 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xoutput310 _1784_/X vssd1 vssd1 vccd1 vccd1 data_out[142] sky130_fd_sc_hd__buf_12
Xoutput343 _1667_/X vssd1 vssd1 vccd1 vccd1 data_out[25] sky130_fd_sc_hd__buf_12
Xoutput321 _1794_/X vssd1 vssd1 vccd1 vccd1 data_out[152] sky130_fd_sc_hd__buf_12
Xoutput332 _1804_/X vssd1 vssd1 vccd1 vccd1 data_out[162] sky130_fd_sc_hd__buf_12
XANTENNA__1166__S _1188_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xoutput365 _1687_/X vssd1 vssd1 vccd1 vccd1 data_out[45] sky130_fd_sc_hd__buf_12
Xoutput354 _1677_/X vssd1 vssd1 vccd1 vccd1 data_out[35] sky130_fd_sc_hd__buf_12
Xoutput387 _1707_/X vssd1 vssd1 vccd1 vccd1 data_out[65] sky130_fd_sc_hd__buf_12
Xoutput376 _1697_/X vssd1 vssd1 vccd1 vccd1 data_out[55] sky130_fd_sc_hd__buf_12
XANTENNA__1156__A1 _2086_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xoutput398 _1717_/X vssd1 vssd1 vccd1 vccd1 data_out[75] sky130_fd_sc_hd__buf_12
XANTENNA__1690__A _2118_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_1529_ _1529_/A1 _1529_/A2 _1529_/B1 _2122_/Q hold266/X vssd1 vssd1 vccd1 vccd1 _1529_/X
+ sky130_fd_sc_hd__a221o_1
XANTENNA__1092__A0 _2210_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__2026__A _2026_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__1631__A2 _1637_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_45_281 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__1395__B2 _2180_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__1147__B2 _1146_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xfanout570 _1519_/A2 vssd1 vssd1 vccd1 vccd1 _1463_/B sky130_fd_sc_hd__clkbuf_4
Xfanout592 _1394_/A vssd1 vssd1 vccd1 vccd1 _1415_/A sky130_fd_sc_hd__clkbuf_4
Xfanout581 _1499_/B1 vssd1 vssd1 vccd1 vccd1 _1503_/B1 sky130_fd_sc_hd__clkbuf_8
XANTENNA__1759__B _1792_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XPHY_90 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__1083__B1 _1095_/B1 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_1880_ _2069_/A vssd1 vssd1 vccd1 vccd1 _1880_/Y sky130_fd_sc_hd__inv_2
XANTENNA__1197__D _1197_/D vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_3_315 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__1775__A _2213_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__1386__B2 _2183_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_51_273 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_3_337 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__1138__A1 _2095_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_1314_ input30/X _1197_/D _1527_/B1 _2207_/Q hold197/X vssd1 vssd1 vccd1 vccd1 _1314_/X
+ sky130_fd_sc_hd__a221o_1
X_2294_ _2312_/CLK _2294_/D _2033_/Y vssd1 vssd1 vccd1 vccd1 _2294_/Q sky130_fd_sc_hd__dfrtp_1
X_1245_ input55/X _1463_/B _1499_/B1 _2230_/Q hold379/X vssd1 vssd1 vccd1 vccd1 _1245_/X
+ sky130_fd_sc_hd__a221o_1
X_1176_ _2168_/Q _2076_/Q _1178_/S vssd1 vssd1 vccd1 vccd1 _1176_/X sky130_fd_sc_hd__mux2_1
XFILLER_0_47_557 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_19_237 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__1074__A0 _2219_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_22 hold178/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_11 hold218/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__1613__A2 _1637_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_27_281 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__1685__A _2113_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_42_251 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__1377__B2 _2186_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__1129__B2 _1128_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_30_457 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_38_557 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__1065__B1 _1095_/B1 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__1368__B2 _2189_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_hold984_A _2165_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_33_262 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_33_284 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_608 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_619 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__1534__S hold80/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_17_12 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__1540__A1 _2116_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_17_45 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_1030_ _2241_/Q hold788/X _1094_/S vssd1 vssd1 vccd1 vccd1 _1030_/X sky130_fd_sc_hd__mux2_1
XFILLER_0_33_33 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_1932_ _1954_/A vssd1 vssd1 vccd1 vccd1 _1932_/Y sky130_fd_sc_hd__inv_2
XFILLER_0_44_549 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_16_229 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_1863_ _1941_/A vssd1 vssd1 vccd1 vccd1 _1863_/Y sky130_fd_sc_hd__inv_2
Xinput31 data_in[127] vssd1 vssd1 vccd1 vccd1 input31/X sky130_fd_sc_hd__buf_1
Xinput20 data_in[117] vssd1 vssd1 vccd1 vccd1 input20/X sky130_fd_sc_hd__clkbuf_1
Xinput53 data_in[147] vssd1 vssd1 vccd1 vccd1 input53/X sky130_fd_sc_hd__clkbuf_2
Xinput42 data_in[137] vssd1 vssd1 vccd1 vccd1 input42/X sky130_fd_sc_hd__clkbuf_1
Xinput64 data_in[157] vssd1 vssd1 vccd1 vccd1 input64/X sky130_fd_sc_hd__buf_1
XANTENNA__1359__B2 _2192_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_1794_ _2232_/Q _1802_/B vssd1 vssd1 vccd1 vccd1 _1794_/X sky130_fd_sc_hd__and2_1
Xinput97 data_in[3] vssd1 vssd1 vccd1 vccd1 input97/X sky130_fd_sc_hd__buf_1
Xinput86 data_in[2] vssd1 vssd1 vccd1 vccd1 input86/X sky130_fd_sc_hd__buf_1
Xinput75 data_in[1] vssd1 vssd1 vccd1 vccd1 input75/X sky130_fd_sc_hd__buf_1
XFILLER_0_12_424 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
Xhold804 la_data_in[2] vssd1 vssd1 vccd1 vccd1 hold15/A sky130_fd_sc_hd__dlygate4sd3_1
Xhold837 _2297_/Q vssd1 vssd1 vccd1 vccd1 hold837/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold815 _2322_/Q vssd1 vssd1 vccd1 vccd1 hold815/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold826 _2253_/Q vssd1 vssd1 vccd1 vccd1 hold826/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold859 _2274_/Q vssd1 vssd1 vccd1 vccd1 hold859/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold848 _2312_/Q vssd1 vssd1 vccd1 vccd1 hold848/X sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA__1444__S hold27/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__1531__B2 _2121_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_2277_ _2291_/CLK _2277_/D _2016_/Y vssd1 vssd1 vccd1 vccd1 _2277_/Q sky130_fd_sc_hd__dfrtp_1
X_1228_ _1227_/X _2235_/Q _1252_/S vssd1 vssd1 vccd1 vccd1 _1228_/X sky130_fd_sc_hd__mux2_1
XFILLER_0_28_3 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_1159_ hold606/X _1189_/A2 _1189_/B1 _1158_/X vssd1 vssd1 vccd1 vccd1 _2265_/D sky130_fd_sc_hd__a22o_1
XFILLER_0_50_508 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA_clkbuf_leaf_23_wb_clk_i_A clkbuf_1_1__f_wb_clk_i/X vssd1 vssd1 vccd1 vccd1
+ sky130_fd_sc_hd__diode_2
XFILLER_0_43_582 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_30_298 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__1522__A1 _2125_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_38_365 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__1589__B2 _2092_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_53_368 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_34_571 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_21_276 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_405 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__1772__B _1792_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__1264__S hold26/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_416 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_427 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_438 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_449 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_2200_ _2212_/CLK _2200_/D _1940_/Y vssd1 vssd1 vccd1 vccd1 _2200_/Q sky130_fd_sc_hd__dfrtp_4
XANTENNA__1513__A1 _1513_/A1 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_2131_ _2223_/CLK _2131_/D _1874_/Y vssd1 vssd1 vccd1 vccd1 _2131_/Q sky130_fd_sc_hd__dfrtp_2
XANTENNA__1513__B2 _2130_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_2062_ _2069_/A vssd1 vssd1 vccd1 vccd1 _2062_/Y sky130_fd_sc_hd__inv_2
X_1013_ _1014_/C _0997_/X _1012_/X _1197_/C _0995_/X vssd1 vssd1 vccd1 vccd1 _1013_/X
+ sky130_fd_sc_hd__a2111o_1
XFILLER_0_17_505 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XANTENNA_clkbuf_1_0__f_wb_clk_i_A clkbuf_0_wb_clk_i/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_1915_ _1916_/A vssd1 vssd1 vccd1 vccd1 _1915_/Y sky130_fd_sc_hd__inv_2
XFILLER_0_44_346 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_1846_ _1916_/A vssd1 vssd1 vccd1 vccd1 _1846_/Y sky130_fd_sc_hd__inv_2
XFILLER_0_4_421 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_13_700 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_13_711 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_1777_ _2215_/Q _1798_/B vssd1 vssd1 vccd1 vccd1 _1777_/X sky130_fd_sc_hd__and2_1
Xhold601 _1137_/X vssd1 vssd1 vccd1 vccd1 _2276_/D sky130_fd_sc_hd__dlygate4sd3_1
Xhold612 hold731/X vssd1 vssd1 vccd1 vccd1 hold612/X sky130_fd_sc_hd__buf_1
XFILLER_0_25_593 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__1963__A _2002_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xhold634 _1067_/X vssd1 vssd1 vccd1 vccd1 _2311_/D sky130_fd_sc_hd__dlygate4sd3_1
Xhold645 hold669/X vssd1 vssd1 vccd1 vccd1 hold645/X sky130_fd_sc_hd__dlymetal6s2s_1
Xhold623 hold691/X vssd1 vssd1 vccd1 vccd1 hold623/X sky130_fd_sc_hd__dlymetal6s2s_1
XANTENNA__1682__B _1715_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xhold667 hold903/X vssd1 vssd1 vccd1 vccd1 hold667/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold656 hold680/X vssd1 vssd1 vccd1 vccd1 hold656/X sky130_fd_sc_hd__buf_1
Xhold678 hold800/X vssd1 vssd1 vccd1 vccd1 hold678/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold689 hold814/X vssd1 vssd1 vccd1 vccd1 hold689/X sky130_fd_sc_hd__dlygate4sd3_1
X_2329_ _2330_/CLK _2329_/D _2068_/Y vssd1 vssd1 vccd1 vccd1 _2329_/Q sky130_fd_sc_hd__dfrtp_1
XFILLER_0_35_335 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_50_305 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__2034__A _2034_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__1440__B1 _1545_/B1 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_16_571 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_16_582 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__1873__A _2002_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_31_585 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XANTENNA_hold947_A _2190_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xinput210 hold264/X vssd1 vssd1 vccd1 vccd1 hold265/A sky130_fd_sc_hd__buf_1
Xinput232 hold382/X vssd1 vssd1 vccd1 vccd1 hold383/A sky130_fd_sc_hd__clkbuf_1
Xinput243 hold5/X vssd1 vssd1 vccd1 vccd1 hold6/A sky130_fd_sc_hd__clkbuf_1
Xinput254 hold551/X vssd1 vssd1 vccd1 vccd1 hold552/A sky130_fd_sc_hd__clkbuf_1
Xinput221 hold371/X vssd1 vssd1 vccd1 vccd1 hold372/A sky130_fd_sc_hd__clkbuf_1
X_1700_ _2128_/Q _1715_/B vssd1 vssd1 vccd1 vccd1 _1700_/X sky130_fd_sc_hd__and2_1
XANTENNA__1431__B1 _1569_/B1 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_53_187 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_41_349 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_1631_ input1/X _1637_/B _1635_/C _2071_/Q hold49/X vssd1 vssd1 vccd1 vccd1 hold50/A
+ sky130_fd_sc_hd__a221o_1
XFILLER_0_30_89 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__1783__A _2221_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_34_390 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_1562_ hold370/X hold987/X hold81/X vssd1 vssd1 vccd1 vccd1 _2105_/D sky130_fd_sc_hd__mux2_1
XTAP_213 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_224 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_202 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_1493_ _1493_/A1 _1503_/A2 _1503_/B1 _2140_/Q hold436/X vssd1 vssd1 vccd1 vccd1 _1493_/X
+ sky130_fd_sc_hd__a221o_1
XFILLER_0_39_65 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_257 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_246 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_235 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_39_98 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_279 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_268 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_55_53 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_2114_ _2173_/CLK _2114_/D _1857_/Y vssd1 vssd1 vccd1 vccd1 _2114_/Q sky130_fd_sc_hd__dfrtp_4
XFILLER_0_55_86 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_2045_ _2065_/A vssd1 vssd1 vccd1 vccd1 _2045_/Y sky130_fd_sc_hd__inv_2
XANTENNA__1958__A _2002_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_29_162 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_32_305 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__1422__B1 _1569_/B1 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_32_327 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_1829_ _1852_/A vssd1 vssd1 vccd1 vccd1 _1829_/Y sky130_fd_sc_hd__inv_2
Xhold420 hold446/X vssd1 vssd1 vccd1 vccd1 hold420/X sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA__1693__A _2121_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xhold453 _1520_/X vssd1 vssd1 vccd1 vccd1 _2126_/D sky130_fd_sc_hd__dlygate4sd3_1
Xhold431 hold563/X vssd1 vssd1 vccd1 vccd1 _1022_/B sky130_fd_sc_hd__buf_1
Xhold442 hold442/A vssd1 vssd1 vccd1 vccd1 _1223_/B sky130_fd_sc_hd__dlygate4sd3_1
Xhold464 _1513_/X vssd1 vssd1 vccd1 vccd1 hold464/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold486 _1453_/X vssd1 vssd1 vccd1 vccd1 _1455_/C sky130_fd_sc_hd__dlygate4sd3_1
Xhold475 _1256_/X vssd1 vssd1 vccd1 vccd1 hold475/X sky130_fd_sc_hd__clkdlybuf4s25_1
Xhold497 la_data_in[61] vssd1 vssd1 vccd1 vccd1 hold497/X sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA__1489__B1 _1503_/B1 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_791 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_780 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__1413__B1 _1545_/B1 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_36_677 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_35_198 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_31_371 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_31_393 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__1542__S hold80/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_output402_A _1721_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_25_78 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_46_408 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__1778__A _2216_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_46_419 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_39_471 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_0993_ hold21/X _1002_/A _1014_/C _0993_/D vssd1 vssd1 vccd1 vccd1 _0993_/X sky130_fd_sc_hd__and4bb_1
XFILLER_0_54_474 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_42_603 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_26_165 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__1404__B1 _1569_/B1 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_42_625 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_14_316 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
Xoutput514 hold590/X vssd1 vssd1 vccd1 vccd1 la_data_out[99] sky130_fd_sc_hd__buf_12
Xoutput503 hold632/X vssd1 vssd1 vccd1 vccd1 la_data_out[88] sky130_fd_sc_hd__buf_12
X_1614_ hold102/X _2079_/Q _1632_/S vssd1 vssd1 vccd1 vccd1 _1614_/X sky130_fd_sc_hd__mux2_1
X_1545_ _1545_/A1 _1198_/A _1545_/B1 _2114_/Q hold44/X vssd1 vssd1 vccd1 vccd1 _1545_/X
+ sky130_fd_sc_hd__a221o_1
XANTENNA__1183__A2 _1183_/A2 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_1476_ hold232/X _2148_/Q _1504_/S vssd1 vssd1 vccd1 vccd1 _1476_/X sky130_fd_sc_hd__mux2_1
XFILLER_0_10_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_2028_ _2033_/A vssd1 vssd1 vccd1 vccd1 _2028_/Y sky130_fd_sc_hd__inv_2
XFILLER_0_49_235 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__1688__A _2116_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_49_279 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_9_343 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_18_600 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_37_419 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_57_290 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_17_110 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_18_633 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA_fanout600_A _1922_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_45_485 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_18_699 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_32_157 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
Xhold250 _1369_/X vssd1 vssd1 vccd1 vccd1 _2188_/D sky130_fd_sc_hd__dlygate4sd3_1
Xhold261 hold261/A vssd1 vssd1 vccd1 vccd1 hold261/X sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_13_393 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_40_190 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xhold283 hold292/X vssd1 vssd1 vccd1 vccd1 hold283/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold294 la_data_in[4] vssd1 vssd1 vccd1 vccd1 hold294/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold272 _1206_/X vssd1 vssd1 vccd1 vccd1 hold272/X sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_51_411 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_23_113 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_24_625 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_23_135 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XANTENNA__1165__A2 _1183_/A2 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_1330_ hold255/X hold961/X hold27/X vssd1 vssd1 vccd1 vccd1 _2201_/D sky130_fd_sc_hd__mux2_1
X_1261_ _1260_/X _2224_/Q hold26/X vssd1 vssd1 vccd1 vccd1 _1261_/X sky130_fd_sc_hd__mux2_1
Xinput7 data_in[105] vssd1 vssd1 vccd1 vccd1 input7/X sky130_fd_sc_hd__buf_1
X_1192_ hold554/X _1192_/B _1192_/C vssd1 vssd1 vccd1 vccd1 _1192_/X sky130_fd_sc_hd__and3b_1
XFILLER_0_36_66 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_52_32 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_46_205 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_46_238 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__1301__A _1310_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_6_324 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XANTENNA__1389__C1 _1388_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_0976_ hold35/X _0977_/B _0977_/C _0976_/D vssd1 vssd1 vccd1 vccd1 _1012_/D sky130_fd_sc_hd__and4_1
XFILLER_0_15_647 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__1447__S hold27/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xoutput300 _1775_/X vssd1 vssd1 vccd1 vccd1 data_out[133] sky130_fd_sc_hd__buf_12
XFILLER_0_42_477 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_42_466 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
Xoutput333 _1658_/X vssd1 vssd1 vccd1 vccd1 data_out[16] sky130_fd_sc_hd__buf_12
Xoutput344 _1668_/X vssd1 vssd1 vccd1 vccd1 data_out[26] sky130_fd_sc_hd__buf_12
Xoutput311 _1785_/X vssd1 vssd1 vccd1 vccd1 data_out[143] sky130_fd_sc_hd__buf_12
Xoutput322 _1795_/X vssd1 vssd1 vccd1 vccd1 data_out[153] sky130_fd_sc_hd__buf_12
XFILLER_0_58_3 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
Xoutput377 _1698_/X vssd1 vssd1 vccd1 vccd1 data_out[56] sky130_fd_sc_hd__buf_12
Xoutput355 _1678_/X vssd1 vssd1 vccd1 vccd1 data_out[36] sky130_fd_sc_hd__buf_12
Xoutput366 _1688_/X vssd1 vssd1 vccd1 vccd1 data_out[46] sky130_fd_sc_hd__buf_12
XANTENNA__1971__A _1979_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xoutput388 _1708_/X vssd1 vssd1 vccd1 vccd1 data_out[66] sky130_fd_sc_hd__buf_12
Xoutput399 _1718_/X vssd1 vssd1 vccd1 vccd1 data_out[76] sky130_fd_sc_hd__buf_12
X_1528_ _1527_/X _2122_/Q hold80/X vssd1 vssd1 vccd1 vccd1 _1528_/X sky130_fd_sc_hd__mux2_1
XANTENNA__1690__B _1724_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_1459_ _1455_/B _0971_/X _1001_/X hold110/X _1810_/C vssd1 vssd1 vccd1 vccd1 _1459_/Y
+ sky130_fd_sc_hd__a41oi_1
XANTENNA__1182__S _1188_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout550_A _1792_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__1092__A1 _2118_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_18_474 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_33_422 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__1395__A2 _1569_/A2 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__2042__A _2065_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_21_617 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_33_477 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_20_127 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__1147__A2 _1189_/A2 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__1881__A _1979_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xfanout560 _1003_/Y vssd1 vssd1 vccd1 vccd1 _1198_/A sky130_fd_sc_hd__clkbuf_4
XANTENNA__1092__S _1188_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xfanout571 _1003_/Y vssd1 vssd1 vccd1 vccd1 _1519_/A2 sky130_fd_sc_hd__buf_4
Xfanout593 _1394_/A vssd1 vssd1 vccd1 vccd1 _1349_/A sky130_fd_sc_hd__clkbuf_2
Xfanout582 _1499_/B1 vssd1 vssd1 vccd1 vccd1 _1495_/B1 sky130_fd_sc_hd__buf_2
XFILLER_0_28_205 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__1607__B1 _1623_/B1 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XPHY_91 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_80 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__1267__S hold26/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_2293_ _2312_/CLK _2293_/D _2032_/Y vssd1 vssd1 vccd1 vccd1 _2293_/Q sky130_fd_sc_hd__dfrtp_1
X_1313_ _1349_/A _1313_/B vssd1 vssd1 vccd1 vccd1 _1313_/X sky130_fd_sc_hd__and2_1
X_1244_ _1271_/A _1244_/B vssd1 vssd1 vccd1 vccd1 _1244_/X sky130_fd_sc_hd__and2_1
X_1175_ hold623/X _1189_/A2 _1189_/B1 _1174_/X vssd1 vssd1 vccd1 vccd1 _2257_/D sky130_fd_sc_hd__a22o_1
XFILLER_0_59_341 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xclkbuf_leaf_19_wb_clk_i clkbuf_1_1__f_wb_clk_i/X vssd1 vssd1 vccd1 vccd1 _2330_/CLK
+ sky130_fd_sc_hd__clkbuf_16
XANTENNA__1074__A1 _2127_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_12 hold135/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_23 hold206/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_35_709 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__1966__A _2039_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_7_666 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_15_411 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__1685__B _1725_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_clkbuf_leaf_13_wb_clk_i_A clkbuf_1_1__f_wb_clk_i/X vssd1 vssd1 vccd1 vccd1
+ sky130_fd_sc_hd__diode_2
X_0959_ hold76/X hold21/X _1002_/A vssd1 vssd1 vccd1 vccd1 _0959_/Y sky130_fd_sc_hd__nor3_1
XANTENNA__1129__A2 _1189_/A2 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout598_A _1913_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_30_469 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__2037__A _2065_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_38_514 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__1876__A _2002_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__1368__A2 _1529_/A2 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_hold977_A _2169_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_21_447 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_609 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_17_57 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_29_514 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_29_547 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_1931_ _1957_/A vssd1 vssd1 vccd1 vccd1 _1931_/Y sky130_fd_sc_hd__inv_2
XFILLER_0_17_709 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__1786__A _2224_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_44_539 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_44_528 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_44_517 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_1862_ _1941_/A vssd1 vssd1 vccd1 vccd1 _1862_/Y sky130_fd_sc_hd__inv_2
Xinput21 data_in[118] vssd1 vssd1 vccd1 vccd1 input21/X sky130_fd_sc_hd__buf_1
Xinput10 data_in[108] vssd1 vssd1 vccd1 vccd1 input10/X sky130_fd_sc_hd__clkbuf_1
Xinput32 data_in[128] vssd1 vssd1 vccd1 vccd1 input32/X sky130_fd_sc_hd__buf_1
Xinput54 data_in[148] vssd1 vssd1 vccd1 vccd1 input54/X sky130_fd_sc_hd__clkbuf_2
Xinput43 data_in[138] vssd1 vssd1 vccd1 vccd1 input43/X sky130_fd_sc_hd__clkbuf_1
XANTENNA__1359__A2 _1529_/A2 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_24_241 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_1793_ _2231_/Q _1804_/B vssd1 vssd1 vccd1 vccd1 _1793_/X sky130_fd_sc_hd__and2_1
Xinput65 data_in[158] vssd1 vssd1 vccd1 vccd1 input65/X sky130_fd_sc_hd__clkbuf_2
Xinput98 data_in[40] vssd1 vssd1 vccd1 vccd1 input98/X sky130_fd_sc_hd__buf_1
Xinput87 data_in[30] vssd1 vssd1 vccd1 vccd1 input87/X sky130_fd_sc_hd__clkbuf_1
Xinput76 data_in[20] vssd1 vssd1 vccd1 vccd1 input76/X sky130_fd_sc_hd__clkbuf_1
XFILLER_0_12_436 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xhold805 _2284_/Q vssd1 vssd1 vccd1 vccd1 hold805/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold827 _2313_/Q vssd1 vssd1 vccd1 vccd1 hold827/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold816 _2254_/Q vssd1 vssd1 vccd1 vccd1 hold816/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold838 _2255_/Q vssd1 vssd1 vccd1 vccd1 hold838/X sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_12_447 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xhold849 _2323_/Q vssd1 vssd1 vccd1 vccd1 hold849/X sky130_fd_sc_hd__dlygate4sd3_1
X_2276_ _2291_/CLK _2276_/D _2015_/Y vssd1 vssd1 vccd1 vccd1 _2276_/Q sky130_fd_sc_hd__dfrtp_1
X_1227_ input62/X _1503_/A2 _1503_/B1 _2236_/Q hold422/X vssd1 vssd1 vccd1 vccd1 _1227_/X
+ sky130_fd_sc_hd__a221o_1
X_1158_ _2177_/Q _2085_/Q _1178_/S vssd1 vssd1 vccd1 vccd1 _1158_/X sky130_fd_sc_hd__mux2_1
XFILLER_0_59_160 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_1089_ hold580/X _1097_/A2 _1097_/B1 _1088_/X vssd1 vssd1 vccd1 vccd1 _2300_/D sky130_fd_sc_hd__a22o_1
XFILLER_0_35_517 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_30_200 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__1589__A2 _1623_/A2 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_53_303 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_53_347 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_34_583 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_21_255 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_21_266 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_406 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_417 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_428 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_439 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__1513__A2 _1519_/A2 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_2130_ _2223_/CLK _2130_/D _1873_/Y vssd1 vssd1 vccd1 vccd1 _2130_/Q sky130_fd_sc_hd__dfrtp_2
X_2061_ _2061_/A vssd1 vssd1 vccd1 vccd1 _2061_/Y sky130_fd_sc_hd__inv_2
X_1012_ _1011_/X _1012_/B _1012_/C _1012_/D vssd1 vssd1 vccd1 vccd1 _1012_/X sky130_fd_sc_hd__and4b_1
XFILLER_0_48_108 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_44_88 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_29_333 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_17_517 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_1914_ _1916_/A vssd1 vssd1 vccd1 vccd1 _1914_/Y sky130_fd_sc_hd__inv_2
X_1845_ _1916_/A vssd1 vssd1 vccd1 vccd1 _1845_/Y sky130_fd_sc_hd__inv_2
XFILLER_0_44_358 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_25_561 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_1776_ _2214_/Q _1802_/B vssd1 vssd1 vccd1 vccd1 _1776_/X sky130_fd_sc_hd__and2_1
Xhold602 hold675/X vssd1 vssd1 vccd1 vccd1 hold602/X sky130_fd_sc_hd__dlymetal6s2s_1
XFILLER_0_12_233 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
Xhold613 _1129_/X vssd1 vssd1 vccd1 vccd1 _2280_/D sky130_fd_sc_hd__dlygate4sd3_1
Xhold635 hold706/X vssd1 vssd1 vccd1 vccd1 hold635/X sky130_fd_sc_hd__buf_1
Xhold624 hold694/X vssd1 vssd1 vccd1 vccd1 hold624/X sky130_fd_sc_hd__dlymetal6s2s_1
XFILLER_0_40_542 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
Xhold668 hold808/X vssd1 vssd1 vccd1 vccd1 hold668/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold657 _1083_/X vssd1 vssd1 vccd1 vccd1 _2303_/D sky130_fd_sc_hd__dlygate4sd3_1
Xhold679 hold807/X vssd1 vssd1 vccd1 vccd1 hold679/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold646 hold713/X vssd1 vssd1 vccd1 vccd1 hold646/X sky130_fd_sc_hd__clkbuf_2
XFILLER_0_40_586 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_40_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_2328_ _2328_/CLK _2328_/D _2067_/Y vssd1 vssd1 vccd1 vccd1 _2328_/Q sky130_fd_sc_hd__dfrtp_1
X_2259_ _2269_/CLK _2259_/D _1998_/Y vssd1 vssd1 vccd1 vccd1 _2259_/Q sky130_fd_sc_hd__dfrtp_1
XFILLER_0_47_141 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_35_325 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__1440__B2 _2165_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_50_317 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__2050__A _2065_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_31_597 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
Xinput200 hold70/X vssd1 vssd1 vccd1 vccd1 hold71/A sky130_fd_sc_hd__clkbuf_1
Xinput211 hold283/X vssd1 vssd1 vccd1 vccd1 hold284/A sky130_fd_sc_hd__clkbuf_1
Xinput222 hold305/X vssd1 vssd1 vccd1 vccd1 hold306/A sky130_fd_sc_hd__clkbuf_1
Xinput244 hold34/X vssd1 vssd1 vccd1 vccd1 hold35/A sky130_fd_sc_hd__clkbuf_1
Xinput233 hold346/X vssd1 vssd1 vccd1 vccd1 hold347/A sky130_fd_sc_hd__buf_1
Xinput255 hold758/X vssd1 vssd1 vccd1 vccd1 _1014_/B sky130_fd_sc_hd__dlymetal6s2s_1
XFILLER_0_14_14 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_39_642 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_39_653 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_53_100 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__1431__B2 _2168_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_1630_ hold32/X _2071_/Q _1632_/S vssd1 vssd1 vccd1 vccd1 hold33/A sky130_fd_sc_hd__mux2_1
XFILLER_0_22_553 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_1561_ input92/X _1623_/A2 _1623_/B1 _2106_/Q hold369/X vssd1 vssd1 vccd1 vccd1 _1561_/X
+ sky130_fd_sc_hd__a221o_1
XANTENNA__1195__A0 hold38/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_1492_ hold411/X _2140_/Q _1520_/S vssd1 vssd1 vccd1 vccd1 _1492_/X sky130_fd_sc_hd__mux2_1
XTAP_214 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_203 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_22_597 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_39_44 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_247 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_236 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_225 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_269 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_258 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_2113_ _2164_/CLK _2113_/D _1856_/Y vssd1 vssd1 vccd1 vccd1 _2113_/Q sky130_fd_sc_hd__dfrtp_4
XANTENNA__1304__A _1310_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_2044_ _2065_/A vssd1 vssd1 vccd1 vccd1 _2044_/Y sky130_fd_sc_hd__inv_2
XANTENNA__1023__B _1811_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_45_612 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_45_623 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_44_100 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_44_166 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_17_358 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__1422__B2 _2171_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_1828_ _1852_/A vssd1 vssd1 vccd1 vccd1 _1828_/Y sky130_fd_sc_hd__inv_2
XANTENNA__1974__A _1979_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_25_380 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xhold410 _1235_/X vssd1 vssd1 vccd1 vccd1 hold410/X sky130_fd_sc_hd__buf_1
XANTENNA__1693__B _1715_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_1759_ _2197_/Q _1792_/B vssd1 vssd1 vccd1 vccd1 _1759_/X sky130_fd_sc_hd__and2_1
Xhold432 _1462_/X vssd1 vssd1 vccd1 vccd1 _1464_/S sky130_fd_sc_hd__dlygate4sd3_1
Xhold454 la_data_in[69] vssd1 vssd1 vccd1 vccd1 hold454/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold421 hold421/A vssd1 vssd1 vccd1 vccd1 _1226_/B sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA__1186__A0 _2163_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xhold443 _1223_/X vssd1 vssd1 vccd1 vccd1 hold443/X sky130_fd_sc_hd__dlymetal6s2s_1
Xhold465 _1514_/X vssd1 vssd1 vccd1 vccd1 _2129_/D sky130_fd_sc_hd__dlygate4sd3_1
Xhold476 _1505_/X vssd1 vssd1 vccd1 vccd1 hold476/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold487 _1455_/X vssd1 vssd1 vccd1 vccd1 hold487/X sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_40_394 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
Xhold498 hold505/X vssd1 vssd1 vccd1 vccd1 hold498/X sky130_fd_sc_hd__clkdlybuf4s25_1
XANTENNA_fanout580_A _1201_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_770 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__1489__A1 _1489_/A1 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_792 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_781 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__1110__A0 _2201_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__2045__A _2065_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_35_111 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_36_623 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_36_645 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__1413__B2 _2174_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__1884__A _2039_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_hold792_A _2116_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__1177__B1 _1183_/B1 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_25_57 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_58_247 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_0992_ _0992_/A _0992_/B hold76/X _1014_/B vssd1 vssd1 vccd1 vccd1 _1012_/B sky130_fd_sc_hd__and4_1
XFILLER_0_39_483 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__1404__B2 _2177_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_41_89 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_14_328 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_2_701 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_41_136 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
Xoutput504 hold636/X vssd1 vssd1 vccd1 vccd1 la_data_out[89] sky130_fd_sc_hd__buf_12
Xoutput515 _2161_/Q vssd1 vssd1 vccd1 vccd1 load_data sky130_fd_sc_hd__buf_12
X_1613_ _1613_/A1 _1637_/B _1635_/C _2080_/Q hold101/X vssd1 vssd1 vccd1 vccd1 _1613_/X
+ sky130_fd_sc_hd__a221o_1
XFILLER_0_41_169 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_1544_ _1543_/X _2114_/Q hold80/X vssd1 vssd1 vccd1 vccd1 _1544_/X sky130_fd_sc_hd__mux2_1
X_1475_ _1475_/A1 _1463_/B _1499_/B1 _2149_/Q hold231/X vssd1 vssd1 vccd1 vccd1 _1475_/X
+ sky130_fd_sc_hd__a221o_1
XFILLER_0_49_214 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_2027_ _2034_/A vssd1 vssd1 vccd1 vccd1 _2027_/Y sky130_fd_sc_hd__inv_2
XFILLER_0_49_225 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_9_300 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__1688__B _1724_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_45_420 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_9_355 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_18_656 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_13_361 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__1159__B1 _1189_/B1 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xhold262 la_data_in[27] vssd1 vssd1 vccd1 vccd1 hold262/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold251 la_data_in[26] vssd1 vssd1 vccd1 vccd1 hold251/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold240 la_data_in[78] vssd1 vssd1 vccd1 vccd1 hold240/X sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_13_372 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xhold284 hold284/A vssd1 vssd1 vccd1 vccd1 _1289_/B sky130_fd_sc_hd__dlygate4sd3_1
Xhold295 hold886/X vssd1 vssd1 vccd1 vccd1 hold295/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold273 _1207_/X vssd1 vssd1 vccd1 vccd1 _2242_/D sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA__1879__A _2065_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__1398__B1 _1529_/B1 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_23_103 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_24_637 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_36_475 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_36_486 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_51_445 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_23_147 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_23_169 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_1260_ input50/X _1519_/A2 _1519_/B1 _2225_/Q hold307/X vssd1 vssd1 vccd1 vccd1 _1260_/X
+ sky130_fd_sc_hd__a221o_1
Xinput8 data_in[106] vssd1 vssd1 vccd1 vccd1 input8/X sky130_fd_sc_hd__buf_1
X_1191_ hold38/X _1191_/B _1191_/C vssd1 vssd1 vccd1 vccd1 _1191_/X sky130_fd_sc_hd__or3_1
XFILLER_0_36_78 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_52_66 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XANTENNA__1625__B2 _2074_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__1389__B1 _1569_/B1 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_0975_ _0971_/C _0969_/C hold561/X _1455_/A vssd1 vssd1 vccd1 vccd1 _0975_/Y sky130_fd_sc_hd__o211ai_1
XFILLER_0_6_336 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_15_615 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_15_626 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_15_659 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xoutput301 _1776_/X vssd1 vssd1 vccd1 vccd1 data_out[134] sky130_fd_sc_hd__buf_12
XFILLER_0_23_670 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
Xoutput334 _1659_/X vssd1 vssd1 vccd1 vccd1 data_out[17] sky130_fd_sc_hd__buf_12
Xoutput312 _1786_/X vssd1 vssd1 vccd1 vccd1 data_out[144] sky130_fd_sc_hd__buf_12
Xoutput323 _1796_/X vssd1 vssd1 vccd1 vccd1 data_out[154] sky130_fd_sc_hd__buf_12
Xoutput345 _1669_/X vssd1 vssd1 vccd1 vccd1 data_out[27] sky130_fd_sc_hd__buf_12
Xoutput367 _1689_/X vssd1 vssd1 vccd1 vccd1 data_out[47] sky130_fd_sc_hd__buf_12
Xoutput356 _1679_/X vssd1 vssd1 vccd1 vccd1 data_out[37] sky130_fd_sc_hd__buf_12
Xoutput378 _1699_/X vssd1 vssd1 vccd1 vccd1 data_out[57] sky130_fd_sc_hd__buf_12
XFILLER_0_10_342 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_2_586 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_22_191 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
Xoutput389 _1709_/X vssd1 vssd1 vccd1 vccd1 data_out[67] sky130_fd_sc_hd__buf_12
XANTENNA__1561__B1 _1623_/B1 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_1527_ _1527_/A1 _1527_/A2 _1527_/B1 _2123_/Q hold285/X vssd1 vssd1 vccd1 vccd1 _1527_/X
+ sky130_fd_sc_hd__a221o_1
X_1458_ hold488/X _2158_/Q _1461_/S vssd1 vssd1 vccd1 vccd1 _1458_/X sky130_fd_sc_hd__mux2_1
X_1389_ input3/X _1569_/A2 _1569_/B1 _2182_/Q _1388_/X vssd1 vssd1 vccd1 vccd1 _1389_/X
+ sky130_fd_sc_hd__a221o_1
XANTENNA__1699__A _2127_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout543_A _1724_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_37_228 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_52_209 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_45_294 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_5_391 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xfanout550 _1792_/B vssd1 vssd1 vccd1 vccd1 _1802_/B sky130_fd_sc_hd__clkbuf_4
Xfanout572 _1201_/X vssd1 vssd1 vccd1 vccd1 _1635_/C sky130_fd_sc_hd__buf_4
Xfanout583 _1519_/B1 vssd1 vssd1 vccd1 vccd1 _1499_/B1 sky130_fd_sc_hd__clkbuf_4
Xfanout561 _1569_/A2 vssd1 vssd1 vccd1 vccd1 _1623_/A2 sky130_fd_sc_hd__buf_4
XANTENNA_hold922_A _2179_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xfanout594 _0952_/Y vssd1 vssd1 vccd1 vccd1 _1394_/A sky130_fd_sc_hd__buf_2
XANTENNA__1607__B2 _2083_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XPHY_92 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__1083__A2 _1095_/A2 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_28_217 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XPHY_70 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_81 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_36_261 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_51_264 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_3_328 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__1543__B1 _1545_/B1 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_47_55 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_2292_ _2312_/CLK _2292_/D _2031_/Y vssd1 vssd1 vccd1 vccd1 _2292_/Q sky130_fd_sc_hd__dfrtp_1
X_1312_ hold13/X _2207_/Q _1318_/S vssd1 vssd1 vccd1 vccd1 hold14/A sky130_fd_sc_hd__mux2_1
X_1243_ hold360/X _2230_/Q _1252_/S vssd1 vssd1 vccd1 vccd1 _1243_/X sky130_fd_sc_hd__mux2_1
X_1174_ _2169_/Q _2077_/Q _1178_/S vssd1 vssd1 vccd1 vccd1 _1174_/X sky130_fd_sc_hd__mux2_1
XFILLER_0_2_57 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_47_548 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_7_612 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA_13 hold256/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_7_645 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA_24 la_data_in[25] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_27_261 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_12_80 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_0958_ _2248_/Q _1445_/A vssd1 vssd1 vccd1 vccd1 _1810_/C sky130_fd_sc_hd__nand2_4
XFILLER_0_27_294 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_42_253 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA_clkbuf_leaf_9_wb_clk_i_A clkbuf_leaf_9_wb_clk_i/A vssd1 vssd1 vccd1 vccd1
+ sky130_fd_sc_hd__diode_2
XANTENNA__1065__A2 _1095_/A2 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_46_570 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__2053__A _2065_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_33_242 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_21_426 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_21_437 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__1525__B1 _1527_/B1 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_33_57 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_1930_ _1941_/A vssd1 vssd1 vccd1 vccd1 _1930_/Y sky130_fd_sc_hd__inv_2
X_1861_ _1941_/A vssd1 vssd1 vccd1 vccd1 _1861_/Y sky130_fd_sc_hd__inv_2
Xinput22 data_in[119] vssd1 vssd1 vccd1 vccd1 input22/X sky130_fd_sc_hd__buf_1
Xinput11 data_in[109] vssd1 vssd1 vccd1 vccd1 input11/X sky130_fd_sc_hd__clkbuf_1
Xinput55 data_in[149] vssd1 vssd1 vccd1 vccd1 input55/X sky130_fd_sc_hd__clkbuf_2
Xinput33 data_in[129] vssd1 vssd1 vccd1 vccd1 input33/X sky130_fd_sc_hd__buf_1
Xinput44 data_in[139] vssd1 vssd1 vccd1 vccd1 input44/X sky130_fd_sc_hd__buf_1
XFILLER_0_24_253 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_1792_ _2230_/Q _1792_/B vssd1 vssd1 vccd1 vccd1 _1792_/X sky130_fd_sc_hd__and2_1
Xinput88 data_in[31] vssd1 vssd1 vccd1 vccd1 input88/X sky130_fd_sc_hd__clkbuf_1
Xinput77 data_in[21] vssd1 vssd1 vccd1 vccd1 input77/X sky130_fd_sc_hd__clkbuf_1
Xinput66 data_in[159] vssd1 vssd1 vccd1 vccd1 input66/X sky130_fd_sc_hd__clkbuf_2
XFILLER_0_3_169 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xhold806 _2269_/Q vssd1 vssd1 vccd1 vccd1 hold806/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold817 _2310_/Q vssd1 vssd1 vccd1 vccd1 hold817/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold828 _2309_/Q vssd1 vssd1 vccd1 vccd1 hold828/X sky130_fd_sc_hd__dlygate4sd3_1
Xinput99 data_in[41] vssd1 vssd1 vccd1 vccd1 input99/X sky130_fd_sc_hd__buf_1
Xhold839 _2265_/Q vssd1 vssd1 vccd1 vccd1 hold839/X sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA__1307__A _1310_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_2275_ _2291_/CLK _2275_/D _2014_/Y vssd1 vssd1 vccd1 vccd1 _2275_/Q sky130_fd_sc_hd__dfrtp_1
X_1226_ _1277_/A _1226_/B vssd1 vssd1 vccd1 vccd1 _1226_/X sky130_fd_sc_hd__and2_1
X_1157_ hold567/X _1157_/A2 _1157_/B1 _1156_/X vssd1 vssd1 vccd1 vccd1 _2266_/D sky130_fd_sc_hd__a22o_1
XFILLER_0_47_312 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_1088_ _2212_/Q _2120_/Q _1112_/S vssd1 vssd1 vccd1 vccd1 _1088_/X sky130_fd_sc_hd__mux2_1
XANTENNA__1977__A _1979_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__1696__B _1715_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__1188__S _1188_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_43_595 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_43_573 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_31_713 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__1507__B1 _1519_/B1 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__1887__A _1979_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_53_315 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_26_518 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_38_378 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_53_337 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_53_326 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_19_581 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__1098__S _1112_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_53_359 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_22_713 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xclkbuf_leaf_4_wb_clk_i clkbuf_leaf_9_wb_clk_i/A vssd1 vssd1 vccd1 vccd1 _2168_/CLK
+ sky130_fd_sc_hd__clkbuf_16
XFILLER_0_21_223 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_407 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_418 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_429 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_28_57 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_2060_ _2069_/A vssd1 vssd1 vccd1 vccd1 _2060_/Y sky130_fd_sc_hd__inv_2
X_1011_ _1002_/A hold21/X vssd1 vssd1 vccd1 vccd1 _1011_/X sky130_fd_sc_hd__and2b_1
XFILLER_0_57_676 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_17_529 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_1913_ _1913_/A vssd1 vssd1 vccd1 vccd1 _1913_/Y sky130_fd_sc_hd__inv_2
XFILLER_0_29_389 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_1844_ _1916_/A vssd1 vssd1 vccd1 vccd1 _1844_/Y sky130_fd_sc_hd__inv_2
XFILLER_0_4_401 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
Xhold603 hold739/X vssd1 vssd1 vccd1 vccd1 hold603/X sky130_fd_sc_hd__clkbuf_2
XFILLER_0_25_573 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_1775_ _2213_/Q _1802_/B vssd1 vssd1 vccd1 vccd1 _1775_/X sky130_fd_sc_hd__and2_1
Xhold636 hold709/X vssd1 vssd1 vccd1 vccd1 hold636/X sky130_fd_sc_hd__dlymetal6s2s_1
Xhold625 hold712/X vssd1 vssd1 vccd1 vccd1 hold625/X sky130_fd_sc_hd__clkbuf_2
Xhold614 hold725/X vssd1 vssd1 vccd1 vccd1 hold614/X sky130_fd_sc_hd__dlymetal6s2s_1
Xhold669 hold863/X vssd1 vssd1 vccd1 vccd1 hold669/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold647 hold716/X vssd1 vssd1 vccd1 vccd1 hold647/X sky130_fd_sc_hd__clkbuf_2
Xhold658 hold672/X vssd1 vssd1 vccd1 vccd1 hold658/X sky130_fd_sc_hd__clkbuf_2
XFILLER_0_40_598 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_2327_ _2328_/CLK _2327_/D _2066_/Y vssd1 vssd1 vccd1 vccd1 _2327_/Q sky130_fd_sc_hd__dfrtp_1
X_2258_ _2296_/CLK _2258_/D _1997_/Y vssd1 vssd1 vccd1 vccd1 _2258_/Q sky130_fd_sc_hd__dfrtp_1
XFILLER_0_33_3 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_1209_ input69/X _1463_/B _1499_/B1 _2242_/Q hold169/X vssd1 vssd1 vccd1 vccd1 _1209_/X
+ sky130_fd_sc_hd__a221o_1
X_2189_ _2194_/CLK _2189_/D _1929_/Y vssd1 vssd1 vccd1 vccd1 _2189_/Q sky130_fd_sc_hd__dfrtp_4
XFILLER_0_48_610 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__1425__C1 hold117/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_47_164 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_35_337 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XANTENNA__1440__A2 _1637_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_43_381 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xinput201 hold42/X vssd1 vssd1 vccd1 vccd1 hold43/A sky130_fd_sc_hd__clkbuf_1
XANTENNA__1381__S _1435_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xinput212 hold351/X vssd1 vssd1 vccd1 vccd1 hold352/A sky130_fd_sc_hd__buf_1
Xinput245 hold490/X vssd1 vssd1 vccd1 vccd1 hold491/A sky130_fd_sc_hd__clkbuf_1
Xinput223 hold473/X vssd1 vssd1 vccd1 vccd1 hold474/A sky130_fd_sc_hd__buf_1
Xinput234 hold420/X vssd1 vssd1 vccd1 vccd1 hold421/A sky130_fd_sc_hd__clkbuf_1
Xinput256 hold75/X vssd1 vssd1 vccd1 vccd1 hold76/A sky130_fd_sc_hd__clkbuf_1
XFILLER_0_39_610 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_39_665 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_39_676 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_53_123 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_26_326 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_38_197 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XANTENNA__1431__A2 _1569_/A2 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_30_25 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_53_167 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__1556__S hold80/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_34_370 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_1560_ hold345/X hold950/X hold81/X vssd1 vssd1 vccd1 vccd1 _2106_/D sky130_fd_sc_hd__mux2_1
X_1491_ _1491_/A1 _1495_/A2 _1495_/B1 _2141_/Q hold410/X vssd1 vssd1 vccd1 vccd1 _1491_/X
+ sky130_fd_sc_hd__a221o_1
XTAP_215 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_204 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_248 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_237 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_226 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_55_11 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__1291__S _1318_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_259 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_2112_ _2164_/CLK _2112_/D _1855_/Y vssd1 vssd1 vccd1 vccd1 _2112_/Q sky130_fd_sc_hd__dfrtp_4
XFILLER_0_12_8 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_2043_ _2065_/A vssd1 vssd1 vccd1 vccd1 _2043_/Y sky130_fd_sc_hd__inv_2
XFILLER_0_17_326 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_17_337 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__1422__A2 _1569_/A2 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_44_178 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_1827_ _1852_/A vssd1 vssd1 vccd1 vccd1 _1827_/Y sky130_fd_sc_hd__inv_2
Xhold411 _1491_/X vssd1 vssd1 vccd1 vccd1 hold411/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold400 hold400/A vssd1 vssd1 vccd1 vccd1 _1283_/B sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA__1466__S _1466_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_1758_ _2196_/Q _1761_/B vssd1 vssd1 vccd1 vccd1 _1758_/X sky130_fd_sc_hd__and2_1
Xhold433 _1464_/X vssd1 vssd1 vccd1 vccd1 _2154_/D sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA__1186__A1 _2071_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_20_80 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
Xhold422 _1226_/X vssd1 vssd1 vccd1 vccd1 hold422/X sky130_fd_sc_hd__clkbuf_2
Xhold444 _1224_/X vssd1 vssd1 vccd1 vccd1 hold444/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold477 _1506_/X vssd1 vssd1 vccd1 vccd1 _2133_/D sky130_fd_sc_hd__dlygate4sd3_1
Xhold466 la_data_in[59] vssd1 vssd1 vccd1 vccd1 hold466/X sky130_fd_sc_hd__dlygate4sd3_1
X_1689_ _2117_/Q _1724_/B vssd1 vssd1 vccd1 vccd1 _1689_/X sky130_fd_sc_hd__and2_1
Xhold455 _1240_/X vssd1 vssd1 vccd1 vccd1 _2231_/D sky130_fd_sc_hd__dlygate4sd3_1
Xhold499 hold499/A vssd1 vssd1 vccd1 vccd1 _1265_/B sky130_fd_sc_hd__dlygate4sd3_1
Xhold488 _1457_/X vssd1 vssd1 vccd1 vccd1 hold488/X sky130_fd_sc_hd__dlygate4sd3_1
XTAP_760 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__1489__A2 _1503_/A2 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_793 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_782 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_771 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_fanout573_A _1201_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__1110__A1 _2109_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_48_473 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_36_635 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_35_156 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_35_189 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_50_137 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__1177__A1 hold658/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_54_410 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_0991_ _0992_/A _0992_/B _1014_/B vssd1 vssd1 vccd1 vccd1 _0991_/X sky130_fd_sc_hd__and3_1
XFILLER_0_41_46 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_41_57 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_26_156 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_27_679 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__1404__A2 _1569_/A2 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_42_616 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_14_307 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_2_713 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_1612_ hold55/X _2080_/Q _1632_/S vssd1 vssd1 vccd1 vccd1 hold56/A sky130_fd_sc_hd__mux2_1
Xoutput505 hold645/X vssd1 vssd1 vccd1 vccd1 la_data_out[90] sky130_fd_sc_hd__buf_12
XFILLER_0_1_223 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xoutput516 _2244_/Q vssd1 vssd1 vccd1 vccd1 load_status[0] sky130_fd_sc_hd__buf_12
XFILLER_0_22_340 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__1168__A1 _2080_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_10_513 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_1543_ _1543_/A1 _1198_/A _1545_/B1 _2115_/Q hold197/X vssd1 vssd1 vccd1 vccd1 _1543_/X
+ sky130_fd_sc_hd__a221o_1
X_1474_ hold170/X _2149_/Q _1504_/S vssd1 vssd1 vccd1 vccd1 _1474_/X sky130_fd_sc_hd__mux2_1
XFILLER_0_5_68 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_5_46 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_2026_ _2026_/A vssd1 vssd1 vccd1 vccd1 _2026_/Y sky130_fd_sc_hd__inv_2
XFILLER_0_49_248 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_9_334 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_45_432 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_32_126 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xhold252 hold295/X vssd1 vssd1 vccd1 vccd1 hold252/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold230 hold230/A vssd1 vssd1 vccd1 vccd1 _1211_/B sky130_fd_sc_hd__dlygate4sd3_1
Xhold241 _1213_/X vssd1 vssd1 vccd1 vccd1 _2240_/D sky130_fd_sc_hd__dlygate4sd3_1
Xhold263 hold263/A vssd1 vssd1 vccd1 vccd1 hold263/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold296 hold303/X vssd1 vssd1 vccd1 vccd1 hold296/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold274 hold278/X vssd1 vssd1 vccd1 vccd1 hold274/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold285 _1289_/X vssd1 vssd1 vccd1 vccd1 hold285/X sky130_fd_sc_hd__buf_1
XTAP_590 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__1619__C1 hold64/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__1095__B1 _1095_/B1 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__2056__A _2069_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_36_421 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XANTENNA__1895__A _2069_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__1398__B2 _2179_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_23_126 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_36_498 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_32_671 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_1190_ _1810_/C hold494/X _2247_/Q vssd1 vssd1 vccd1 vccd1 _1190_/X sky130_fd_sc_hd__o21a_1
Xinput9 data_in[107] vssd1 vssd1 vccd1 vccd1 input9/X sky130_fd_sc_hd__clkbuf_1
XFILLER_0_59_502 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__1086__A0 _2213_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__1625__A2 _1637_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_52_78 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_39_281 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_54_251 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__1389__B2 _2182_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_6_348 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_0974_ _0971_/C hold755/X hold561/X _1455_/A vssd1 vssd1 vccd1 vccd1 _0974_/X sky130_fd_sc_hd__o211a_1
XFILLER_0_42_424 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_15_638 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xoutput335 _1660_/X vssd1 vssd1 vccd1 vccd1 data_out[18] sky130_fd_sc_hd__buf_12
Xoutput313 _1787_/X vssd1 vssd1 vccd1 vccd1 data_out[145] sky130_fd_sc_hd__buf_12
Xoutput302 _1777_/X vssd1 vssd1 vccd1 vccd1 data_out[135] sky130_fd_sc_hd__buf_12
Xoutput324 _1797_/X vssd1 vssd1 vccd1 vccd1 data_out[155] sky130_fd_sc_hd__buf_12
XFILLER_0_2_565 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xoutput368 _1690_/X vssd1 vssd1 vccd1 vccd1 data_out[48] sky130_fd_sc_hd__buf_12
Xoutput357 _1680_/X vssd1 vssd1 vccd1 vccd1 data_out[38] sky130_fd_sc_hd__buf_12
Xoutput346 _1670_/X vssd1 vssd1 vccd1 vccd1 data_out[28] sky130_fd_sc_hd__buf_12
X_1526_ _1525_/X _2123_/Q hold80/X vssd1 vssd1 vccd1 vccd1 _1526_/X sky130_fd_sc_hd__mux2_1
Xoutput379 _1700_/X vssd1 vssd1 vccd1 vccd1 data_out[58] sky130_fd_sc_hd__buf_12
XANTENNA__1561__B2 _2106_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_1457_ _1198_/X _1456_/X hold487/X _1545_/B1 vssd1 vssd1 vccd1 vccd1 _1457_/X sky130_fd_sc_hd__a211o_1
X_1388_ _1394_/A hold2/X vssd1 vssd1 vccd1 vccd1 _1388_/X sky130_fd_sc_hd__and2_2
XANTENNA__1699__B _1715_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__1077__B1 _1095_/B1 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_2009_ _2034_/A vssd1 vssd1 vccd1 vccd1 _2009_/Y sky130_fd_sc_hd__inv_2
XANTENNA_fanout536_A hold80/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_33_457 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xfanout540 _1724_/B vssd1 vssd1 vccd1 vccd1 _1725_/B sky130_fd_sc_hd__clkbuf_4
Xfanout551 _1641_/Y vssd1 vssd1 vccd1 vccd1 _1792_/B sky130_fd_sc_hd__clkbuf_4
Xfanout562 _1569_/A2 vssd1 vssd1 vccd1 vccd1 _1619_/A2 sky130_fd_sc_hd__clkbuf_4
Xfanout584 _1201_/X vssd1 vssd1 vccd1 vccd1 _1519_/B1 sky130_fd_sc_hd__buf_4
Xfanout573 _1201_/X vssd1 vssd1 vccd1 vccd1 _1545_/B1 sky130_fd_sc_hd__clkbuf_4
Xfanout595 _1310_/A vssd1 vssd1 vccd1 vccd1 _1277_/A sky130_fd_sc_hd__buf_2
XANTENNA__1068__A0 _2222_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__1607__A2 _1623_/A2 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_22_15 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XPHY_60 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_71 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_82 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_93 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_24_402 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_36_251 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA_output288_A _1764_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_2291_ _2291_/CLK _2291_/D _2030_/Y vssd1 vssd1 vccd1 vccd1 _2291_/Q sky130_fd_sc_hd__dfrtp_1
XANTENNA__1543__B2 _2115_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_1311_ input31/X _1197_/D _1541_/B1 _2208_/Q hold12/X vssd1 vssd1 vccd1 vccd1 hold13/A
+ sky130_fd_sc_hd__a221o_1
X_1242_ input57/X _1495_/A2 _1495_/B1 _2231_/Q hold359/X vssd1 vssd1 vccd1 vccd1 _1242_/X
+ sky130_fd_sc_hd__a221o_1
X_1173_ hold638/X _1183_/A2 _1183_/B1 _1172_/X vssd1 vssd1 vccd1 vccd1 _2258_/D sky130_fd_sc_hd__a22o_1
XANTENNA__1059__B1 _1097_/B1 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_14 _1191_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_25 hold94/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_0957_ _2248_/Q _1445_/A vssd1 vssd1 vccd1 vccd1 _1455_/A sky130_fd_sc_hd__and2_2
XFILLER_0_15_446 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_30_438 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__1474__S _1504_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_1509_ _1509_/A1 _1519_/A2 _1519_/B1 _2132_/Q hold373/X vssd1 vssd1 vccd1 vccd1 _1509_/X
+ sky130_fd_sc_hd__a221o_1
XFILLER_0_46_560 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_18_251 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_18_262 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_34_711 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_33_221 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_33_254 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__1384__S _1435_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_21_449 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__1525__A1 _1525_/A1 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_17_15 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_29_505 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_1860_ _1949_/A vssd1 vssd1 vccd1 vccd1 _1860_/Y sky130_fd_sc_hd__inv_2
Xinput12 data_in[10] vssd1 vssd1 vccd1 vccd1 input12/X sky130_fd_sc_hd__buf_1
X_1791_ _2229_/Q _1804_/B vssd1 vssd1 vccd1 vccd1 _1791_/X sky130_fd_sc_hd__and2_1
Xinput45 data_in[13] vssd1 vssd1 vccd1 vccd1 input45/X sky130_fd_sc_hd__buf_1
Xinput23 data_in[11] vssd1 vssd1 vccd1 vccd1 input23/X sky130_fd_sc_hd__buf_1
Xinput34 data_in[12] vssd1 vssd1 vccd1 vccd1 input34/X sky130_fd_sc_hd__buf_1
Xinput89 data_in[32] vssd1 vssd1 vccd1 vccd1 input89/X sky130_fd_sc_hd__clkbuf_1
Xinput78 data_in[22] vssd1 vssd1 vccd1 vccd1 input78/X sky130_fd_sc_hd__clkbuf_1
Xinput56 data_in[14] vssd1 vssd1 vccd1 vccd1 input56/X sky130_fd_sc_hd__buf_1
Xinput67 data_in[15] vssd1 vssd1 vccd1 vccd1 input67/X sky130_fd_sc_hd__clkbuf_1
Xhold807 _2315_/Q vssd1 vssd1 vccd1 vccd1 hold807/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold818 _2268_/Q vssd1 vssd1 vccd1 vccd1 hold818/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold829 _2328_/Q vssd1 vssd1 vccd1 vccd1 hold829/X sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA__1294__S _1318_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_58_44 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_2274_ _2291_/CLK _2274_/D _2013_/Y vssd1 vssd1 vccd1 vccd1 _2274_/Q sky130_fd_sc_hd__dfrtp_1
X_1225_ hold444/X _2236_/Q _1252_/S vssd1 vssd1 vccd1 vccd1 _1225_/X sky130_fd_sc_hd__mux2_1
X_1156_ _2178_/Q _2086_/Q _1156_/S vssd1 vssd1 vccd1 vccd1 _1156_/X sky130_fd_sc_hd__mux2_1
X_1087_ _2301_/Q _1095_/A2 _1095_/B1 _1086_/X vssd1 vssd1 vccd1 vccd1 _1087_/X sky130_fd_sc_hd__a22o_1
XFILLER_0_7_432 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_23_80 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_35_508 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_7_465 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_28_582 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_1989_ _2008_/A vssd1 vssd1 vccd1 vccd1 _1989_/Y sky130_fd_sc_hd__inv_2
XFILLER_0_15_221 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_30_246 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__1507__A1 _1507_/A1 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_38_324 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XANTENNA__2064__A _2069_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__1443__B1 _1545_/B1 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_19_593 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_34_541 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA_hold982_A _2099_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_21_235 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_21_279 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_408 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_419 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_1010_ _0986_/A _1001_/X _1008_/Y _1009_/X vssd1 vssd1 vccd1 vccd1 _1194_/A sky130_fd_sc_hd__o211ai_1
X_1912_ _1913_/A vssd1 vssd1 vccd1 vccd1 _1912_/Y sky130_fd_sc_hd__inv_2
XFILLER_0_29_379 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__1434__B1 _1569_/B1 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_1843_ _1916_/A vssd1 vssd1 vccd1 vccd1 _1843_/Y sky130_fd_sc_hd__inv_2
XFILLER_0_4_424 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_4_413 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_25_585 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_1774_ _2212_/Q _1804_/B vssd1 vssd1 vccd1 vccd1 _1774_/X sky130_fd_sc_hd__and2_1
XFILLER_0_12_213 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xhold604 hold735/X vssd1 vssd1 vccd1 vccd1 hold604/X sky130_fd_sc_hd__clkbuf_2
Xhold615 hold720/X vssd1 vssd1 vccd1 vccd1 hold615/X sky130_fd_sc_hd__buf_1
Xhold626 hold700/X vssd1 vssd1 vccd1 vccd1 hold626/X sky130_fd_sc_hd__clkbuf_2
XFILLER_0_40_533 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xhold648 hold660/X vssd1 vssd1 vccd1 vccd1 hold648/X sky130_fd_sc_hd__buf_1
Xhold637 hold690/X vssd1 vssd1 vccd1 vccd1 hold637/X sky130_fd_sc_hd__buf_1
Xhold659 hold794/X vssd1 vssd1 vccd1 vccd1 hold659/X sky130_fd_sc_hd__dlygate4sd3_1
X_2326_ _2328_/CLK _2326_/D _2065_/Y vssd1 vssd1 vccd1 vccd1 _2326_/Q sky130_fd_sc_hd__dfrtp_1
X_2257_ _2269_/CLK _2257_/D _1996_/Y vssd1 vssd1 vccd1 vccd1 _2257_/Q sky130_fd_sc_hd__dfrtp_1
X_1208_ _1277_/A _1208_/B vssd1 vssd1 vccd1 vccd1 _1208_/X sky130_fd_sc_hd__and2_1
XFILLER_0_26_3 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_2188_ _2219_/CLK _2188_/D _1928_/Y vssd1 vssd1 vccd1 vccd1 _2188_/Q sky130_fd_sc_hd__dfrtp_4
X_1139_ hold597/X _1139_/A2 _1139_/B1 _1138_/X vssd1 vssd1 vccd1 vccd1 _2275_/D sky130_fd_sc_hd__a22o_1
XFILLER_0_47_110 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__1425__B1 _1569_/B1 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_48_677 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA_fanout616_A _2039_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_35_349 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_43_360 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_7_295 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_43_393 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_31_544 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xinput202 hold195/X vssd1 vssd1 vccd1 vccd1 hold196/A sky130_fd_sc_hd__clkbuf_1
Xinput235 hold441/X vssd1 vssd1 vccd1 vccd1 hold442/A sky130_fd_sc_hd__clkbuf_1
Xinput224 hold315/X vssd1 vssd1 vccd1 vccd1 hold316/A sky130_fd_sc_hd__clkbuf_1
Xinput213 hold399/X vssd1 vssd1 vccd1 vccd1 hold400/A sky130_fd_sc_hd__clkbuf_1
Xinput257 hold108/X vssd1 vssd1 vccd1 vccd1 hold109/A sky130_fd_sc_hd__clkbuf_1
Xinput246 hold558/X vssd1 vssd1 vccd1 vccd1 _0977_/D sky130_fd_sc_hd__dlymetal6s2s_1
XANTENNA__2059__A _2069_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__1898__A _1949_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__1416__B1 _1545_/B1 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_53_113 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_19_390 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_30_15 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_34_360 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_1490_ hold385/X _2141_/Q _1504_/S vssd1 vssd1 vccd1 vccd1 _1490_/X sky130_fd_sc_hd__mux2_1
XTAP_205 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_238 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_216 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_227 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_39_68 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_249 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold1 hold1/A vssd1 vssd1 vccd1 vccd1 hold1/X sky130_fd_sc_hd__dlygate4sd3_1
X_2111_ _2164_/CLK _2111_/D _1854_/Y vssd1 vssd1 vccd1 vccd1 _2111_/Q sky130_fd_sc_hd__dfrtp_4
XANTENNA_clkbuf_leaf_22_wb_clk_i_A clkbuf_1_1__f_wb_clk_i/X vssd1 vssd1 vccd1 vccd1
+ sky130_fd_sc_hd__diode_2
X_2042_ _2065_/A vssd1 vssd1 vccd1 vccd1 _2042_/Y sky130_fd_sc_hd__inv_2
XFILLER_0_29_121 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_57_452 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_45_603 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_9_549 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_29_132 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__1407__B1 _1569_/B1 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_44_135 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_32_319 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_1826_ _1852_/A vssd1 vssd1 vccd1 vccd1 _1826_/Y sky130_fd_sc_hd__inv_2
XFILLER_0_25_393 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
Xhold401 _1283_/X vssd1 vssd1 vccd1 vccd1 hold401/X sky130_fd_sc_hd__buf_1
X_1757_ _2195_/Q _1792_/B vssd1 vssd1 vccd1 vccd1 _1757_/X sky130_fd_sc_hd__and2_1
Xhold423 _1485_/X vssd1 vssd1 vccd1 vccd1 hold423/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold445 _1225_/X vssd1 vssd1 vccd1 vccd1 _2236_/D sky130_fd_sc_hd__dlygate4sd3_1
Xhold412 _1492_/X vssd1 vssd1 vccd1 vccd1 _2140_/D sky130_fd_sc_hd__dlygate4sd3_1
Xhold434 hold454/X vssd1 vssd1 vccd1 vccd1 hold434/X sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_40_341 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XANTENNA__1591__C1 hold521/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xhold467 _1270_/X vssd1 vssd1 vccd1 vccd1 _2221_/D sky130_fd_sc_hd__dlygate4sd3_1
Xhold456 la_data_in[32] vssd1 vssd1 vccd1 vccd1 hold456/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold478 la_data_in[63] vssd1 vssd1 vccd1 vccd1 hold478/X sky130_fd_sc_hd__dlygate4sd3_1
X_1688_ _2116_/Q _1724_/B vssd1 vssd1 vccd1 vccd1 _1688_/X sky130_fd_sc_hd__and2_1
Xhold489 _1458_/X vssd1 vssd1 vccd1 vccd1 _2158_/D sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA__1482__S _1504_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_761 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_750 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_794 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_783 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_772 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_2309_ _2315_/CLK _2309_/D _2048_/Y vssd1 vssd1 vccd1 vccd1 _2309_/Q sky130_fd_sc_hd__dfrtp_1
XFILLER_0_29_90 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA_fanout566_A _1527_/A2 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_48_452 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_0_80 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_35_113 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_36_669 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_50_127 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_31_330 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__1177__A2 _1183_/A2 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_31_374 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xhold990 _2093_/Q vssd1 vssd1 vccd1 vccd1 hold990/X sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA_hold945_A _2127_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_58_227 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_0990_ _0990_/A _1012_/D _1012_/C _0990_/D vssd1 vssd1 vccd1 vccd1 _1197_/C sky130_fd_sc_hd__and4_2
XFILLER_0_42_628 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_1611_ input12/X _1637_/B _1635_/C _2081_/Q hold54/X vssd1 vssd1 vccd1 vccd1 hold55/A
+ sky130_fd_sc_hd__a221o_1
XFILLER_0_50_661 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
Xoutput506 hold575/X vssd1 vssd1 vccd1 vccd1 la_data_out[91] sky130_fd_sc_hd__buf_12
Xoutput517 _2245_/Q vssd1 vssd1 vccd1 vccd1 load_status[1] sky130_fd_sc_hd__buf_12
XANTENNA__1573__C1 hold290/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_1542_ _1541_/X _2115_/Q hold80/X vssd1 vssd1 vccd1 vccd1 _1542_/X sky130_fd_sc_hd__mux2_1
X_1473_ _1473_/A1 _1463_/B _1499_/B1 _2150_/Q hold169/X vssd1 vssd1 vccd1 vccd1 _1473_/X
+ sky130_fd_sc_hd__a221o_1
X_2025_ _2026_/A vssd1 vssd1 vccd1 vccd1 _2025_/Y sky130_fd_sc_hd__inv_2
XFILLER_0_15_92 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_18_603 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_45_444 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_17_124 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_1809_ _1809_/A _1809_/B _1635_/B vssd1 vssd1 vccd1 vccd1 _1810_/D sky130_fd_sc_hd__or3b_1
XANTENNA__1159__A2 _1189_/A2 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xhold220 _1605_/X vssd1 vssd1 vccd1 vccd1 hold220/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold253 hold253/A vssd1 vssd1 vccd1 vccd1 _1328_/B sky130_fd_sc_hd__dlygate4sd3_1
Xhold242 hold260/X vssd1 vssd1 vccd1 vccd1 hold261/A sky130_fd_sc_hd__dlygate4sd3_1
Xhold231 _1211_/X vssd1 vssd1 vccd1 vccd1 hold231/X sky130_fd_sc_hd__buf_1
Xhold286 _1290_/X vssd1 vssd1 vccd1 vccd1 hold286/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold275 hold275/A vssd1 vssd1 vccd1 vccd1 _1355_/B sky130_fd_sc_hd__dlygate4sd3_1
Xhold264 hold319/X vssd1 vssd1 vccd1 vccd1 hold264/X sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_40_193 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
Xhold297 hold297/A vssd1 vssd1 vccd1 vccd1 _1214_/B sky130_fd_sc_hd__dlygate4sd3_1
XTAP_580 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_591 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_36_411 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_36_433 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XANTENNA__1387__S _1435_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_51_414 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__1398__A2 _1529_/A2 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_32_694 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__1086__A1 _2121_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_59_558 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_46_208 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_54_230 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__1389__A2 _1569_/A2 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_0973_ _0977_/C _0973_/B _0973_/C _0973_/D vssd1 vssd1 vccd1 vccd1 _0973_/X sky130_fd_sc_hd__or4_1
XFILLER_0_15_617 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_27_455 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__1297__S _1318_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_30_609 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
Xoutput303 _1778_/X vssd1 vssd1 vccd1 vccd1 data_out[136] sky130_fd_sc_hd__buf_12
Xoutput314 _1788_/X vssd1 vssd1 vccd1 vccd1 data_out[146] sky130_fd_sc_hd__buf_12
Xoutput325 _1798_/X vssd1 vssd1 vccd1 vccd1 data_out[156] sky130_fd_sc_hd__buf_12
Xoutput369 _1691_/X vssd1 vssd1 vccd1 vccd1 data_out[49] sky130_fd_sc_hd__buf_12
Xoutput347 _1671_/X vssd1 vssd1 vccd1 vccd1 data_out[29] sky130_fd_sc_hd__buf_12
Xoutput336 _1661_/X vssd1 vssd1 vccd1 vccd1 data_out[19] sky130_fd_sc_hd__buf_12
Xoutput358 _1681_/X vssd1 vssd1 vccd1 vccd1 data_out[39] sky130_fd_sc_hd__buf_12
X_1525_ _1525_/A1 _1527_/A2 _1527_/B1 _2124_/Q hold353/X vssd1 vssd1 vccd1 vccd1 _1525_/X
+ sky130_fd_sc_hd__a221o_1
XANTENNA__1561__A2 _1623_/A2 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_1456_ hold2/X hold88/X vssd1 vssd1 vccd1 vccd1 _1456_/X sky130_fd_sc_hd__xor2_1
X_1387_ hold522/X hold975/X _1435_/S vssd1 vssd1 vccd1 vccd1 _2182_/D sky130_fd_sc_hd__mux2_1
XANTENNA__1077__B2 _1076_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_2008_ _2008_/A vssd1 vssd1 vccd1 vccd1 _2008_/Y sky130_fd_sc_hd__inv_2
XANTENNA_fanout529_A _1157_/A2 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_18_477 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_33_414 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_21_609 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_5_393 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_14_672 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xfanout541 _1680_/B vssd1 vssd1 vccd1 vccd1 _1677_/B sky130_fd_sc_hd__clkbuf_4
Xfanout530 _1022_/X vssd1 vssd1 vccd1 vccd1 _1157_/A2 sky130_fd_sc_hd__clkbuf_4
Xfanout552 _1157_/B1 vssd1 vssd1 vccd1 vccd1 _1189_/B1 sky130_fd_sc_hd__buf_4
Xfanout563 _1003_/Y vssd1 vssd1 vccd1 vccd1 _1569_/A2 sky130_fd_sc_hd__clkbuf_8
Xfanout574 _1569_/B1 vssd1 vssd1 vccd1 vccd1 _1623_/B1 sky130_fd_sc_hd__buf_4
Xfanout585 _1112_/S vssd1 vssd1 vccd1 vccd1 _1188_/S sky130_fd_sc_hd__clkbuf_8
Xfanout596 _1310_/A vssd1 vssd1 vccd1 vccd1 _1271_/A sky130_fd_sc_hd__clkbuf_2
XANTENNA__2067__A _2069_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__1068__A1 _2130_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XPHY_83 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_50 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_28_208 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XPHY_61 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_72 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_49_591 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XPHY_94 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_22_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_22_49 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_52_701 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_47_46 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_2290_ _2312_/CLK _2290_/D _2029_/Y vssd1 vssd1 vccd1 vccd1 _2290_/Q sky130_fd_sc_hd__dfrtp_1
X_1310_ _1310_/A hold11/X vssd1 vssd1 vccd1 vccd1 hold12/A sky130_fd_sc_hd__and2_1
XFILLER_0_47_68 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_47_57 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_1241_ _1271_/A _1241_/B vssd1 vssd1 vccd1 vccd1 _1241_/X sky130_fd_sc_hd__and2_1
X_1172_ _2170_/Q _2078_/Q _1188_/S vssd1 vssd1 vccd1 vccd1 _1172_/X sky130_fd_sc_hd__mux2_1
XFILLER_0_19_208 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XANTENNA_26 _1415_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_27_252 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA_15 _1358_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_12_71 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_15_414 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_0956_ _1988_/A vssd1 vssd1 vccd1 vccd1 _0956_/Y sky130_fd_sc_hd__inv_2
XFILLER_0_42_233 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_12_93 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_2_341 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_2_363 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_56_3 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_1508_ hold308/X _2132_/Q _1520_/S vssd1 vssd1 vccd1 vccd1 _1508_/X sky130_fd_sc_hd__mux2_1
XANTENNA__1490__S _1504_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_1439_ _1445_/A hold16/X vssd1 vssd1 vccd1 vccd1 hold17/A sky130_fd_sc_hd__and2_1
XANTENNA__1470__A1 _2151_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_18_230 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_34_701 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__1525__A2 _1527_/A2 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_33_15 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_37_561 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
Xinput13 data_in[110] vssd1 vssd1 vccd1 vccd1 input13/X sky130_fd_sc_hd__clkbuf_1
X_1790_ _2228_/Q _1804_/B vssd1 vssd1 vccd1 vccd1 _1790_/X sky130_fd_sc_hd__and2_1
Xinput35 data_in[130] vssd1 vssd1 vccd1 vccd1 input35/X sky130_fd_sc_hd__buf_1
Xinput24 data_in[120] vssd1 vssd1 vccd1 vccd1 input24/X sky130_fd_sc_hd__buf_1
Xinput46 data_in[140] vssd1 vssd1 vccd1 vccd1 input46/X sky130_fd_sc_hd__buf_1
XFILLER_0_24_233 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
Xinput57 data_in[150] vssd1 vssd1 vccd1 vccd1 input57/X sky130_fd_sc_hd__clkbuf_2
Xinput68 data_in[160] vssd1 vssd1 vccd1 vccd1 input68/X sky130_fd_sc_hd__clkbuf_2
Xinput79 data_in[23] vssd1 vssd1 vccd1 vccd1 input79/X sky130_fd_sc_hd__buf_1
XFILLER_0_52_586 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
Xhold808 _2316_/Q vssd1 vssd1 vccd1 vccd1 hold808/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold819 _2270_/Q vssd1 vssd1 vccd1 vccd1 hold819/X sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_12_439 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_20_494 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_2273_ _2291_/CLK _2273_/D _2012_/Y vssd1 vssd1 vccd1 vccd1 _2273_/Q sky130_fd_sc_hd__dfrtp_1
X_1224_ input63/X _1503_/A2 _1503_/B1 _2237_/Q hold443/X vssd1 vssd1 vccd1 vccd1 _1224_/X
+ sky130_fd_sc_hd__a221o_1
X_1155_ hold607/X _1189_/A2 _1189_/B1 _1154_/X vssd1 vssd1 vccd1 vccd1 _2267_/D sky130_fd_sc_hd__a22o_1
X_1086_ _2213_/Q _2121_/Q _1086_/S vssd1 vssd1 vccd1 vccd1 _1086_/X sky130_fd_sc_hd__mux2_1
XFILLER_0_59_141 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_47_369 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_16_701 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_28_561 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_23_92 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_1988_ _1988_/A vssd1 vssd1 vccd1 vccd1 _1988_/Y sky130_fd_sc_hd__inv_2
XFILLER_0_43_586 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_31_704 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA_fanout596_A _1310_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__1507__A2 _1519_/A2 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_3_91 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__1140__A0 _2186_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_38_336 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_53_306 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__1443__B2 _2164_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__1443__A1 _1443_/A1 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_19_561 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_34_520 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_34_531 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA_hold975_A _2182_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_21_225 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_34_597 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_21_247 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_409 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_28_15 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XANTENNA_clkbuf_leaf_12_wb_clk_i_A clkbuf_1_1__f_wb_clk_i/X vssd1 vssd1 vccd1 vccd1
+ sky130_fd_sc_hd__diode_2
X_1911_ _1913_/A vssd1 vssd1 vccd1 vccd1 _1911_/Y sky130_fd_sc_hd__inv_2
XANTENNA__1434__B2 _2167_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_1842_ _1916_/A vssd1 vssd1 vccd1 vccd1 _1842_/Y sky130_fd_sc_hd__inv_2
XFILLER_0_25_542 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_52_361 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_1773_ _2211_/Q _1804_/B vssd1 vssd1 vccd1 vccd1 _1773_/X sky130_fd_sc_hd__and2_1
Xhold605 hold728/X vssd1 vssd1 vccd1 vccd1 hold605/X sky130_fd_sc_hd__dlymetal6s2s_1
XFILLER_0_8_58 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xhold616 hold710/X vssd1 vssd1 vccd1 vccd1 hold616/X sky130_fd_sc_hd__buf_1
Xhold627 hold723/X vssd1 vssd1 vccd1 vccd1 hold627/X sky130_fd_sc_hd__clkbuf_2
XFILLER_0_25_597 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
Xhold638 hold687/X vssd1 vssd1 vccd1 vccd1 hold638/X sky130_fd_sc_hd__clkbuf_2
Xhold649 hold692/X vssd1 vssd1 vccd1 vccd1 hold649/X sky130_fd_sc_hd__clkbuf_2
XFILLER_0_0_642 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_2325_ _2328_/CLK _2325_/D _2064_/Y vssd1 vssd1 vccd1 vccd1 _2325_/Q sky130_fd_sc_hd__dfrtp_1
X_2256_ _2256_/CLK _2256_/D _1995_/Y vssd1 vssd1 vccd1 vccd1 _2256_/Q sky130_fd_sc_hd__dfrtp_1
XANTENNA__1122__A0 _2195_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_1207_ hold272/X _2242_/Q _1252_/S vssd1 vssd1 vccd1 vccd1 _1207_/X sky130_fd_sc_hd__mux2_1
X_2187_ _2219_/CLK _2187_/D _1927_/Y vssd1 vssd1 vccd1 vccd1 _2187_/Q sky130_fd_sc_hd__dfrtp_4
XFILLER_0_19_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_1138_ _2187_/Q _2095_/Q _1156_/S vssd1 vssd1 vccd1 vccd1 _1138_/X sky130_fd_sc_hd__mux2_1
X_1069_ hold576/X _1097_/A2 _1097_/B1 _1068_/X vssd1 vssd1 vccd1 vccd1 _2310_/D sky130_fd_sc_hd__a22o_1
XANTENNA__1425__B2 _2170_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_47_144 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA_fanout609_A _2026_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__1189__B1 _1189_/B1 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_16_586 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_31_512 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xclkbuf_leaf_12_wb_clk_i clkbuf_1_1__f_wb_clk_i/X vssd1 vssd1 vccd1 vccd1 _2224_/CLK
+ sky130_fd_sc_hd__clkbuf_16
Xinput225 hold323/X vssd1 vssd1 vccd1 vccd1 hold324/A sky130_fd_sc_hd__clkbuf_1
Xinput236 hold513/X vssd1 vssd1 vccd1 vccd1 hold514/A sky130_fd_sc_hd__clkbuf_1
Xinput214 hold389/X vssd1 vssd1 vccd1 vccd1 hold390/A sky130_fd_sc_hd__clkbuf_1
Xinput203 hold10/X vssd1 vssd1 vccd1 vccd1 hold11/A sky130_fd_sc_hd__clkbuf_1
Xinput258 hold20/X vssd1 vssd1 vccd1 vccd1 hold21/A sky130_fd_sc_hd__clkbuf_1
Xinput247 hold754/X vssd1 vssd1 vccd1 vccd1 _0977_/C sky130_fd_sc_hd__clkbuf_2
XANTENNA__1113__B1 _1183_/B1 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_39_623 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_39_645 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__1416__B2 _2173_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_39_656 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_53_136 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_53_169 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_53_158 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA_output263_A _1642_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_206 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_239 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_217 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_228 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_55_35 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xhold2 hold2/A vssd1 vssd1 vccd1 vccd1 hold2/X sky130_fd_sc_hd__clkbuf_2
X_2110_ _2164_/CLK _2110_/D _1853_/Y vssd1 vssd1 vccd1 vccd1 _2110_/Q sky130_fd_sc_hd__dfrtp_4
X_2041_ _2061_/A vssd1 vssd1 vccd1 vccd1 _2041_/Y sky130_fd_sc_hd__inv_2
XANTENNA__1104__A0 _2204_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_29_111 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__1407__B2 _2176_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_45_615 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_53_670 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_25_361 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_1825_ _1852_/A vssd1 vssd1 vccd1 vccd1 _1825_/Y sky130_fd_sc_hd__inv_2
XFILLER_0_32_309 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_1756_ _2194_/Q _1756_/B vssd1 vssd1 vccd1 vccd1 _1756_/X sky130_fd_sc_hd__and2_1
Xhold402 _1523_/X vssd1 vssd1 vccd1 vccd1 hold402/X sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_25_383 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xhold435 hold435/A vssd1 vssd1 vccd1 vccd1 _1238_/B sky130_fd_sc_hd__dlygate4sd3_1
Xhold413 hold480/X vssd1 vssd1 vccd1 vccd1 hold413/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold424 la_data_in[80] vssd1 vssd1 vccd1 vccd1 hold424/X sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA__1591__B1 _1623_/B1 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xhold457 la_data_in[19] vssd1 vssd1 vccd1 vccd1 hold1/A sky130_fd_sc_hd__dlygate4sd3_1
Xhold446 la_data_in[73] vssd1 vssd1 vccd1 vccd1 hold446/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold468 hold482/X vssd1 vssd1 vccd1 vccd1 hold468/X sky130_fd_sc_hd__dlygate4sd3_1
X_1687_ _2115_/Q _1724_/B vssd1 vssd1 vccd1 vccd1 _1687_/X sky130_fd_sc_hd__and2_2
Xhold479 _1258_/X vssd1 vssd1 vccd1 vccd1 _2225_/D sky130_fd_sc_hd__dlygate4sd3_1
XTAP_751 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_740 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_784 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_795 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_773 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_762 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_2308_ _2330_/CLK _2308_/D _2047_/Y vssd1 vssd1 vccd1 vccd1 _2308_/Q sky130_fd_sc_hd__dfrtp_1
X_2239_ _2239_/CLK _2239_/D _1979_/Y vssd1 vssd1 vccd1 vccd1 _2239_/Q sky130_fd_sc_hd__dfrtp_1
XANTENNA_fanout559_A _1003_/Y vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_35_103 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_36_615 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_23_309 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_35_169 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xhold980 _2090_/Q vssd1 vssd1 vccd1 vccd1 hold980/X sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_8_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xhold991 _2110_/Q vssd1 vssd1 vccd1 vccd1 hold991/X sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA_hold938_A _2096_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__1702__A _2130_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_27_615 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_41_15 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_26_136 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_39_497 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_14_309 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_1610_ hold157/X _2081_/Q hold80/X vssd1 vssd1 vccd1 vccd1 _1610_/X sky130_fd_sc_hd__mux2_1
Xoutput507 hold576/X vssd1 vssd1 vccd1 vccd1 la_data_out[92] sky130_fd_sc_hd__buf_12
Xoutput518 _2246_/Q vssd1 vssd1 vccd1 vccd1 load_status[2] sky130_fd_sc_hd__buf_12
X_1541_ _1541_/A1 _1197_/D _1541_/B1 _2116_/Q hold12/X vssd1 vssd1 vccd1 vccd1 _1541_/X
+ sky130_fd_sc_hd__a221o_1
X_1472_ _1471_/X _2150_/Q _1504_/S vssd1 vssd1 vccd1 vccd1 _1472_/X sky130_fd_sc_hd__mux2_1
X_2024_ _2033_/A vssd1 vssd1 vccd1 vccd1 _2024_/Y sky130_fd_sc_hd__inv_2
XANTENNA__1628__A1 _2072_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_49_239 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_9_358 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_18_659 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_1808_ hold2/A hold88/A _1808_/C _1808_/D vssd1 vssd1 vccd1 vccd1 _1809_/A sky130_fd_sc_hd__or4_1
Xhold210 hold891/X vssd1 vssd1 vccd1 vccd1 hold210/X sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_13_331 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_13_353 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_1739_ _2177_/Q _1761_/B vssd1 vssd1 vccd1 vccd1 _1739_/X sky130_fd_sc_hd__and2_1
Xhold243 hold243/A vssd1 vssd1 vccd1 vccd1 _1352_/B sky130_fd_sc_hd__dlygate4sd3_1
Xhold221 hold256/X vssd1 vssd1 vccd1 vccd1 hold221/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold232 _1475_/X vssd1 vssd1 vccd1 vccd1 hold232/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold287 _1291_/X vssd1 vssd1 vccd1 vccd1 _2214_/D sky130_fd_sc_hd__dlygate4sd3_1
Xhold265 hold265/A vssd1 vssd1 vccd1 vccd1 _1292_/B sky130_fd_sc_hd__dlygate4sd3_1
Xhold254 _1328_/X vssd1 vssd1 vccd1 vccd1 hold254/X sky130_fd_sc_hd__buf_1
Xhold276 _1355_/X vssd1 vssd1 vccd1 vccd1 hold276/X sky130_fd_sc_hd__dlymetal6s2s_1
Xhold298 _1214_/X vssd1 vssd1 vccd1 vccd1 hold298/X sky130_fd_sc_hd__dlymetal6s2s_1
XTAP_570 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_581 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_592 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__1619__B2 _2077_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__1095__A2 _1095_/A2 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_48_250 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_36_445 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_31_183 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_36_15 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_52_36 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_27_401 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_39_250 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_0972_ _0977_/C _0976_/D _0973_/D vssd1 vssd1 vccd1 vccd1 _0972_/X sky130_fd_sc_hd__or3_1
XFILLER_0_27_445 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_54_264 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_54_297 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_42_448 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xoutput304 _1779_/X vssd1 vssd1 vccd1 vccd1 data_out[137] sky130_fd_sc_hd__buf_12
XFILLER_0_50_470 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xoutput315 _1789_/X vssd1 vssd1 vccd1 vccd1 data_out[147] sky130_fd_sc_hd__buf_12
Xoutput326 _1799_/X vssd1 vssd1 vccd1 vccd1 data_out[157] sky130_fd_sc_hd__buf_12
XFILLER_0_22_161 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
Xoutput359 _1645_/X vssd1 vssd1 vccd1 vccd1 data_out[3] sky130_fd_sc_hd__buf_12
Xoutput348 _1644_/X vssd1 vssd1 vccd1 vccd1 data_out[2] sky130_fd_sc_hd__buf_12
Xoutput337 _1643_/X vssd1 vssd1 vccd1 vccd1 data_out[1] sky130_fd_sc_hd__buf_12
X_1524_ hold402/X _2124_/Q hold80/X vssd1 vssd1 vccd1 vccd1 _1524_/X sky130_fd_sc_hd__mux2_1
XFILLER_0_10_345 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_1455_ _1455_/A _1455_/B _1455_/C _1455_/D vssd1 vssd1 vccd1 vccd1 _1455_/X sky130_fd_sc_hd__and4_1
X_1386_ input4/X _1533_/A2 _1529_/B1 _2183_/Q hold521/X vssd1 vssd1 vccd1 vccd1 _1386_/X
+ sky130_fd_sc_hd__a221o_1
X_2007_ _2026_/A vssd1 vssd1 vccd1 vccd1 _2007_/Y sky130_fd_sc_hd__inv_2
XANTENNA__1077__A2 _1095_/A2 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__1488__S _1504_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_45_297 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_5_361 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_14_662 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_13_183 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__1537__B1 _1541_/B1 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xfanout531 _1097_/A2 vssd1 vssd1 vccd1 vccd1 _1095_/A2 sky130_fd_sc_hd__buf_4
Xfanout542 _1724_/B vssd1 vssd1 vccd1 vccd1 _1680_/B sky130_fd_sc_hd__clkbuf_4
Xfanout575 _1569_/B1 vssd1 vssd1 vccd1 vccd1 _1619_/B1 sky130_fd_sc_hd__clkbuf_4
XANTENNA_hold469_A hold469/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xfanout553 _1157_/B1 vssd1 vssd1 vccd1 vccd1 _1139_/B1 sky130_fd_sc_hd__clkbuf_4
Xfanout564 _1527_/A2 vssd1 vssd1 vccd1 vccd1 _1197_/D sky130_fd_sc_hd__buf_4
Xfanout597 _0952_/Y vssd1 vssd1 vccd1 vccd1 _1310_/A sky130_fd_sc_hd__buf_4
Xfanout586 _1112_/S vssd1 vssd1 vccd1 vccd1 _1178_/S sky130_fd_sc_hd__clkbuf_8
XPHY_40 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_51 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_62 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_73 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_95 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_84 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_52_713 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_36_264 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_51_245 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_20_632 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_20_687 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_1240_ _1239_/X _2231_/Q _1252_/S vssd1 vssd1 vccd1 vccd1 _1240_/X sky130_fd_sc_hd__mux2_1
X_1171_ hold624/X _1189_/A2 _1189_/B1 _1170_/X vssd1 vssd1 vccd1 vccd1 _2259_/D sky130_fd_sc_hd__a22o_1
XANTENNA__1059__A2 _1097_/A2 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_55_551 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA_16 la_data_in[30] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_7_648 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_12_61 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_15_426 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_0955_ _2243_/Q vssd1 vssd1 vccd1 vccd1 _0955_/Y sky130_fd_sc_hd__inv_2
XFILLER_0_42_256 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XANTENNA__1519__B1 _1519_/B1 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_23_481 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_1507_ _1507_/A1 _1519_/A2 _1519_/B1 _2133_/Q hold307/X vssd1 vssd1 vccd1 vccd1 _1507_/X
+ sky130_fd_sc_hd__a221o_1
XFILLER_0_49_3 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_1438_ _1437_/X _2165_/Q hold27/X vssd1 vssd1 vccd1 vccd1 _1438_/X sky130_fd_sc_hd__mux2_1
X_1369_ hold249/X _2188_/Q _1372_/S vssd1 vssd1 vccd1 vccd1 _1369_/X sky130_fd_sc_hd__mux2_1
XFILLER_0_18_242 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_46_573 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_18_297 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_33_267 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_56_326 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_37_551 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_37_573 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
Xinput36 data_in[131] vssd1 vssd1 vccd1 vccd1 input36/X sky130_fd_sc_hd__buf_1
Xinput25 data_in[121] vssd1 vssd1 vccd1 vccd1 input25/X sky130_fd_sc_hd__buf_1
Xinput14 data_in[111] vssd1 vssd1 vccd1 vccd1 input14/X sky130_fd_sc_hd__clkbuf_1
Xinput69 data_in[161] vssd1 vssd1 vccd1 vccd1 input69/X sky130_fd_sc_hd__clkbuf_2
Xinput58 data_in[151] vssd1 vssd1 vccd1 vccd1 input58/X sky130_fd_sc_hd__clkbuf_2
Xinput47 data_in[141] vssd1 vssd1 vccd1 vccd1 input47/X sky130_fd_sc_hd__buf_1
Xhold809 _2300_/Q vssd1 vssd1 vccd1 vccd1 hold809/X sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_20_473 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_2272_ _2291_/CLK _2272_/D _2011_/Y vssd1 vssd1 vccd1 vccd1 _2272_/Q sky130_fd_sc_hd__dfrtp_1
X_1223_ _1277_/A _1223_/B vssd1 vssd1 vccd1 vccd1 _1223_/X sky130_fd_sc_hd__and2_1
X_1154_ _2179_/Q _2087_/Q _1178_/S vssd1 vssd1 vccd1 vccd1 _1154_/X sky130_fd_sc_hd__mux2_1
X_1085_ hold652/X _1095_/A2 _1095_/B1 _1084_/X vssd1 vssd1 vccd1 vccd1 _2302_/D sky130_fd_sc_hd__a22o_1
XFILLER_0_47_304 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_47_337 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_1987_ _1988_/A vssd1 vssd1 vccd1 vccd1 _1987_/Y sky130_fd_sc_hd__inv_2
XFILLER_0_16_713 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_43_532 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_43_576 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_43_598 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA_fanout589_A _1094_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__1140__A1 _2094_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__1428__C1 hold64/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_19_551 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_38_348 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_53_329 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_19_573 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_34_510 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_34_587 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA_hold968_A _2199_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_28_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_44_15 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_57_613 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA_clkbuf_leaf_8_wb_clk_i_A clkbuf_leaf_9_wb_clk_i/A vssd1 vssd1 vccd1 vccd1
+ sky130_fd_sc_hd__diode_2
XFILLER_0_29_337 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_1910_ _1916_/A vssd1 vssd1 vccd1 vccd1 _1910_/Y sky130_fd_sc_hd__inv_2
XANTENNA__1434__A2 _1569_/A2 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_1841_ _1922_/A vssd1 vssd1 vccd1 vccd1 _1841_/Y sky130_fd_sc_hd__inv_2
XFILLER_0_25_532 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_1772_ _2210_/Q _1792_/B vssd1 vssd1 vccd1 vccd1 _1772_/X sky130_fd_sc_hd__and2_1
XFILLER_0_52_373 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
Xhold617 hold718/X vssd1 vssd1 vccd1 vccd1 hold617/X sky130_fd_sc_hd__dlymetal6s2s_1
Xhold606 hold740/X vssd1 vssd1 vccd1 vccd1 hold606/X sky130_fd_sc_hd__clkbuf_2
XFILLER_0_40_524 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
Xhold628 hold729/X vssd1 vssd1 vccd1 vccd1 hold628/X sky130_fd_sc_hd__clkbuf_2
Xhold639 hold711/X vssd1 vssd1 vccd1 vccd1 hold639/X sky130_fd_sc_hd__clkbuf_2
X_2324_ _2330_/CLK _2324_/D _2063_/Y vssd1 vssd1 vccd1 vccd1 _2324_/Q sky130_fd_sc_hd__dfrtp_1
X_2255_ _2291_/CLK _2255_/D _1994_/Y vssd1 vssd1 vccd1 vccd1 _2255_/Q sky130_fd_sc_hd__dfrtp_1
X_1206_ input70/X _1197_/D hold271/X vssd1 vssd1 vccd1 vccd1 _1206_/X sky130_fd_sc_hd__a21o_1
X_2186_ _2212_/CLK _2186_/D _1926_/Y vssd1 vssd1 vccd1 vccd1 _2186_/Q sky130_fd_sc_hd__dfrtp_4
XANTENNA__1122__A1 _2103_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_1137_ _2276_/Q _1139_/A2 _1139_/B1 _1136_/X vssd1 vssd1 vccd1 vccd1 _1137_/X sky130_fd_sc_hd__a22o_1
X_1068_ _2222_/Q _2130_/Q _1086_/S vssd1 vssd1 vccd1 vccd1 _1068_/X sky130_fd_sc_hd__mux2_1
XANTENNA__1425__A2 _1569_/A2 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_47_123 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_47_167 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_16_510 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_35_329 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_16_521 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__1496__S _1504_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_16_565 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_43_384 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_11_270 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
Xinput226 hold310/X vssd1 vssd1 vccd1 vccd1 hold311/A sky130_fd_sc_hd__clkbuf_1
Xinput215 hold448/X vssd1 vssd1 vccd1 vccd1 hold449/A sky130_fd_sc_hd__clkbuf_1
Xinput204 hold57/X vssd1 vssd1 vccd1 vccd1 hold58/A sky130_fd_sc_hd__clkbuf_1
Xinput237 hold413/X vssd1 vssd1 vccd1 vccd1 hold414/A sky130_fd_sc_hd__clkbuf_1
Xinput248 hold539/X vssd1 vssd1 vccd1 vccd1 hold540/A sky130_fd_sc_hd__buf_1
Xinput259 hold99/X vssd1 vssd1 vccd1 vccd1 hold100/A sky130_fd_sc_hd__clkbuf_1
XFILLER_0_14_29 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_39_613 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__1416__A2 _1637_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_39_668 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_39_679 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_26_329 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_38_189 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_19_381 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_34_373 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_39_15 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_218 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_229 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_207 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold3 hold3/A vssd1 vssd1 vccd1 vccd1 hold3/X sky130_fd_sc_hd__dlygate4sd3_1
X_2040_ _2065_/A vssd1 vssd1 vccd1 vccd1 _2040_/Y sky130_fd_sc_hd__inv_2
XANTENNA__1104__A1 _2112_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__1407__A2 _1003_/Y vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_5_713 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_1824_ _1988_/A vssd1 vssd1 vccd1 vccd1 _1824_/Y sky130_fd_sc_hd__inv_2
X_1755_ _2193_/Q _1756_/B vssd1 vssd1 vccd1 vccd1 _1755_/X sky130_fd_sc_hd__and2_1
XFILLER_0_25_373 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
Xhold403 _1524_/X vssd1 vssd1 vccd1 vccd1 _2124_/D sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_52_192 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_52_181 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xhold414 hold414/A vssd1 vssd1 vccd1 vccd1 _1217_/B sky130_fd_sc_hd__dlygate4sd3_1
Xhold425 _1472_/X vssd1 vssd1 vccd1 vccd1 _2150_/D sky130_fd_sc_hd__dlygate4sd3_1
Xhold436 _1238_/X vssd1 vssd1 vccd1 vccd1 hold436/X sky130_fd_sc_hd__buf_1
XANTENNA__1591__B2 _2091_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xhold447 _1228_/X vssd1 vssd1 vccd1 vccd1 _2235_/D sky130_fd_sc_hd__dlygate4sd3_1
Xhold458 hold1/X vssd1 vssd1 vccd1 vccd1 hold458/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold469 hold469/A vssd1 vssd1 vccd1 vccd1 _1271_/B sky130_fd_sc_hd__dlygate4sd3_1
X_1686_ _2114_/Q _1725_/B vssd1 vssd1 vccd1 vccd1 _1686_/X sky130_fd_sc_hd__and2_1
XTAP_752 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_741 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_730 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_785 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_774 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_763 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_2307_ _2328_/CLK _2307_/D _2046_/Y vssd1 vssd1 vccd1 vccd1 _2307_/Q sky130_fd_sc_hd__dfrtp_1
X_2238_ _2238_/CLK _2238_/D _1978_/Y vssd1 vssd1 vccd1 vccd1 _2238_/Q sky130_fd_sc_hd__dfrtp_1
XTAP_796 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_31_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_2169_ _2182_/CLK _2169_/D _1909_/Y vssd1 vssd1 vccd1 vccd1 _2169_/Q sky130_fd_sc_hd__dfrtp_4
XFILLER_0_45_91 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_48_421 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_48_443 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_48_432 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_36_605 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_36_627 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_35_159 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_16_362 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_43_181 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_31_387 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
Xhold981 _2092_/Q vssd1 vssd1 vccd1 vccd1 hold981/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold970 _2180_/Q vssd1 vssd1 vccd1 vccd1 hold970/X sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_31_398 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xhold992 _2173_/Q vssd1 vssd1 vccd1 vccd1 hold992/X sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA__1702__B _1715_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__1098__A0 _2207_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_39_410 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_35_671 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xoutput508 hold633/X vssd1 vssd1 vccd1 vccd1 la_data_out[93] sky130_fd_sc_hd__buf_12
XFILLER_0_22_321 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_1540_ _1539_/X _2116_/Q hold80/X vssd1 vssd1 vccd1 vccd1 _1540_/X sky130_fd_sc_hd__mux2_1
XANTENNA__1573__B2 _2100_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xoutput519 _2155_/Q vssd1 vssd1 vccd1 vccd1 master_ena_proc sky130_fd_sc_hd__buf_12
XFILLER_0_22_365 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_1471_ _1471_/A1 _1197_/D _1541_/B1 _2151_/Q hold271/X vssd1 vssd1 vccd1 vccd1 _1471_/X
+ sky130_fd_sc_hd__a221o_1
X_2023_ _2033_/A vssd1 vssd1 vccd1 vccd1 _2023_/Y sky130_fd_sc_hd__inv_2
XANTENNA__1104__S _1188_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__1089__B1 _1097_/B1 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_45_402 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_17_104 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_45_479 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_1807_ _1807_/A _1807_/B vssd1 vssd1 vccd1 vccd1 _2243_/D sky130_fd_sc_hd__nor2_1
XFILLER_0_31_82 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_32_129 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
Xhold211 la_data_in[25] vssd1 vssd1 vccd1 vccd1 hold211/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold200 _1540_/X vssd1 vssd1 vccd1 vccd1 _2116_/D sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_25_192 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
Xhold222 hold222/A vssd1 vssd1 vccd1 vccd1 _1361_/B sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_13_376 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
Xhold233 _1476_/X vssd1 vssd1 vccd1 vccd1 _2148_/D sky130_fd_sc_hd__dlygate4sd3_1
Xhold244 _1352_/X vssd1 vssd1 vccd1 vccd1 hold244/X sky130_fd_sc_hd__dlymetal6s2s_1
X_1738_ _2176_/Q _1761_/B vssd1 vssd1 vccd1 vccd1 _1738_/X sky130_fd_sc_hd__and2_1
Xhold277 _1356_/X vssd1 vssd1 vccd1 vccd1 hold277/X sky130_fd_sc_hd__dlygate4sd3_1
X_1669_ _2097_/Q _1677_/B vssd1 vssd1 vccd1 vccd1 _1669_/X sky130_fd_sc_hd__and2_1
Xhold266 _1292_/X vssd1 vssd1 vccd1 vccd1 hold266/X sky130_fd_sc_hd__buf_1
Xhold255 _1329_/X vssd1 vssd1 vccd1 vccd1 hold255/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold299 _1477_/X vssd1 vssd1 vccd1 vccd1 hold299/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold288 hold301/X vssd1 vssd1 vccd1 vccd1 hold288/X sky130_fd_sc_hd__dlygate4sd3_1
XTAP_560 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_fanout571_A _1003_/Y vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_571 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_582 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_593 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_48_262 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_51_405 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_8_381 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_23_129 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_51_449 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_31_162 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__1555__B2 _2109_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_hold950_A _2106_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_36_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_59_505 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_52_15 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_52_48 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_39_262 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_6_307 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_0971_ _0978_/A _0978_/B _0971_/C _0970_/X vssd1 vssd1 vccd1 vccd1 _0971_/X sky130_fd_sc_hd__or4b_1
XFILLER_0_15_608 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_42_427 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_50_460 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xoutput305 _1780_/X vssd1 vssd1 vccd1 vccd1 data_out[138] sky130_fd_sc_hd__buf_12
Xoutput316 _1790_/X vssd1 vssd1 vccd1 vccd1 data_out[148] sky130_fd_sc_hd__buf_12
Xoutput338 _1662_/X vssd1 vssd1 vccd1 vccd1 data_out[20] sky130_fd_sc_hd__buf_12
Xoutput349 _1672_/X vssd1 vssd1 vccd1 vccd1 data_out[30] sky130_fd_sc_hd__buf_12
X_1523_ _1523_/A1 _1527_/A2 _1527_/B1 _2125_/Q hold401/X vssd1 vssd1 vccd1 vccd1 _1523_/X
+ sky130_fd_sc_hd__a221o_1
XFILLER_0_50_493 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xoutput327 _1800_/X vssd1 vssd1 vccd1 vccd1 data_out[158] sky130_fd_sc_hd__buf_12
X_1454_ _0953_/Y _0990_/A _1014_/C hold22/X vssd1 vssd1 vccd1 vccd1 _1455_/D sky130_fd_sc_hd__a31oi_1
X_1385_ _1394_/A _1385_/B vssd1 vssd1 vccd1 vccd1 _1385_/X sky130_fd_sc_hd__and2_1
X_2006_ _2008_/A vssd1 vssd1 vccd1 vccd1 _2006_/Y sky130_fd_sc_hd__inv_2
XFILLER_0_26_82 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_33_427 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_33_438 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_5_373 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XANTENNA__1537__A1 _1537_/A1 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__1537__B2 _2118_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xfanout532 _1097_/A2 vssd1 vssd1 vccd1 vccd1 _1057_/A2 sky130_fd_sc_hd__clkbuf_4
Xfanout521 hold26/X vssd1 vssd1 vccd1 vccd1 hold27/A sky130_fd_sc_hd__clkbuf_1
Xfanout554 _1157_/B1 vssd1 vssd1 vccd1 vccd1 _1183_/B1 sky130_fd_sc_hd__buf_4
Xfanout565 _1529_/A2 vssd1 vssd1 vccd1 vccd1 _1533_/A2 sky130_fd_sc_hd__buf_4
Xfanout543 _1724_/B vssd1 vssd1 vccd1 vccd1 _1715_/B sky130_fd_sc_hd__clkbuf_4
Xfanout587 _1112_/S vssd1 vssd1 vccd1 vccd1 _1156_/S sky130_fd_sc_hd__buf_4
Xfanout598 _1913_/A vssd1 vssd1 vccd1 vccd1 _1988_/A sky130_fd_sc_hd__buf_8
XTAP_390 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xfanout576 _1201_/X vssd1 vssd1 vccd1 vccd1 _1569_/B1 sky130_fd_sc_hd__clkbuf_8
XPHY_30 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_41 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_52 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_63 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_74 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_37_700 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XPHY_96 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_85 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_22_29 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_24_405 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_51_279 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xclkbuf_leaf_7_wb_clk_i clkbuf_leaf_9_wb_clk_i/A vssd1 vssd1 vccd1 vccd1 _2217_/CLK
+ sky130_fd_sc_hd__clkbuf_16
XFILLER_0_20_699 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_1170_ _2171_/Q _2079_/Q _1188_/S vssd1 vssd1 vccd1 vccd1 _1170_/X sky130_fd_sc_hd__mux2_1
XFILLER_0_47_508 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA_17 la_data_in[34] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_42_213 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_0954_ _1025_/B vssd1 vssd1 vccd1 vccd1 _1810_/B sky130_fd_sc_hd__inv_2
XFILLER_0_15_405 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_15_438 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_15_449 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_42_268 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_23_460 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__1519__B2 _2127_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__1519__A1 _1519_/A1 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_2_365 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_1506_ hold476/X _2133_/Q _1520_/S vssd1 vssd1 vccd1 vccd1 _1506_/X sky130_fd_sc_hd__mux2_1
X_1437_ _1437_/A1 _1198_/A _1545_/B1 _2166_/Q hold176/X vssd1 vssd1 vccd1 vccd1 _1437_/X
+ sky130_fd_sc_hd__a221o_1
X_1368_ input10/X _1529_/A2 _1533_/B1 _2189_/Q hold248/X vssd1 vssd1 vccd1 vccd1 _1368_/X
+ sky130_fd_sc_hd__a221o_1
X_1299_ input36/X _1529_/A2 _1529_/B1 _2212_/Q hold147/X vssd1 vssd1 vccd1 vccd1 _1299_/X
+ sky130_fd_sc_hd__a221o_1
XANTENNA_fanout534_A hold80/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_38_519 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_33_279 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__1446__B1 _1545_/B1 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_29_508 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_37_585 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
Xinput26 data_in[122] vssd1 vssd1 vccd1 vccd1 input26/X sky130_fd_sc_hd__buf_1
Xinput15 data_in[112] vssd1 vssd1 vccd1 vccd1 input15/X sky130_fd_sc_hd__clkbuf_1
Xinput37 data_in[132] vssd1 vssd1 vccd1 vccd1 input37/X sky130_fd_sc_hd__buf_1
Xinput59 data_in[152] vssd1 vssd1 vccd1 vccd1 input59/X sky130_fd_sc_hd__clkbuf_2
Xinput48 data_in[142] vssd1 vssd1 vccd1 vccd1 input48/X sky130_fd_sc_hd__buf_1
XFILLER_0_12_419 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_24_246 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA_output453_A hold658/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_2271_ _2291_/CLK _2271_/D _2010_/Y vssd1 vssd1 vccd1 vccd1 _2271_/Q sky130_fd_sc_hd__dfrtp_1
X_1222_ _1221_/X _2237_/Q _1252_/S vssd1 vssd1 vccd1 vccd1 _1222_/X sky130_fd_sc_hd__mux2_1
XANTENNA__1901__A _1949_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_1153_ hold570/X _1157_/A2 _1157_/B1 _1152_/X vssd1 vssd1 vccd1 vccd1 _2268_/D sky130_fd_sc_hd__a22o_1
X_1084_ _2214_/Q _2122_/Q _1086_/S vssd1 vssd1 vccd1 vccd1 _1084_/X sky130_fd_sc_hd__mux2_1
XANTENNA__1437__B1 _1545_/B1 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__1112__S _1112_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_47_349 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_7_424 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_1986_ _1988_/A vssd1 vssd1 vccd1 vccd1 _1986_/Y sky130_fd_sc_hd__inv_2
XFILLER_0_7_468 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_43_566 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_43_555 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_15_279 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__1811__A _1811_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__1428__B1 _1569_/B1 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_19_585 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_19_596 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_34_533 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_21_216 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__1705__B _1724_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_28_39 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_44_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__1419__B1 _1545_/B1 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_29_349 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_1840_ _1922_/A vssd1 vssd1 vccd1 vccd1 _1840_/Y sky130_fd_sc_hd__inv_2
XFILLER_0_37_393 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_1771_ _2209_/Q _1804_/B vssd1 vssd1 vccd1 vccd1 _1771_/X sky130_fd_sc_hd__and2_1
Xhold618 hold705/X vssd1 vssd1 vccd1 vccd1 hold618/X sky130_fd_sc_hd__dlymetal6s2s_1
Xhold607 hold738/X vssd1 vssd1 vccd1 vccd1 hold607/X sky130_fd_sc_hd__clkbuf_2
XFILLER_0_40_536 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xhold629 hold722/X vssd1 vssd1 vccd1 vccd1 hold629/X sky130_fd_sc_hd__clkbuf_2
X_2323_ _2330_/CLK _2323_/D _2062_/Y vssd1 vssd1 vccd1 vccd1 _2323_/Q sky130_fd_sc_hd__dfrtp_1
XFILLER_0_0_699 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_18_50 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_2254_ _2269_/CLK _2254_/D _1993_/Y vssd1 vssd1 vccd1 vccd1 _2254_/Q sky130_fd_sc_hd__dfrtp_1
X_1205_ _1277_/A _1205_/B vssd1 vssd1 vccd1 vccd1 _1205_/X sky130_fd_sc_hd__and2_1
X_2185_ _2212_/CLK _2185_/D _1925_/Y vssd1 vssd1 vccd1 vccd1 _2185_/Q sky130_fd_sc_hd__dfrtp_4
X_1136_ _2188_/Q _2096_/Q _1156_/S vssd1 vssd1 vccd1 vccd1 _1136_/X sky130_fd_sc_hd__mux2_1
XFILLER_0_47_113 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_1067_ _2311_/Q _1095_/A2 _1095_/B1 _1066_/X vssd1 vssd1 vccd1 vccd1 _1067_/X sky130_fd_sc_hd__a22o_1
XFILLER_0_34_71 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_47_135 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_34_93 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_16_533 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__1189__A2 _1189_/A2 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_1969_ _1982_/A vssd1 vssd1 vccd1 vccd1 _1969_/Y sky130_fd_sc_hd__inv_2
XFILLER_0_31_503 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_31_547 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_31_558 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
Xinput227 hold377/X vssd1 vssd1 vccd1 vccd1 hold378/A sky130_fd_sc_hd__clkbuf_1
Xinput205 hold93/X vssd1 vssd1 vccd1 vccd1 hold94/A sky130_fd_sc_hd__clkbuf_1
Xinput216 hold338/X vssd1 vssd1 vccd1 vccd1 hold339/A sky130_fd_sc_hd__buf_1
Xinput238 hold296/X vssd1 vssd1 vccd1 vccd1 hold297/A sky130_fd_sc_hd__clkbuf_1
Xinput249 hold484/X vssd1 vssd1 vccd1 vccd1 _0979_/A sky130_fd_sc_hd__buf_1
XANTENNA__1113__A2 _1183_/A2 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xclkbuf_leaf_21_wb_clk_i clkbuf_1_1__f_wb_clk_i/X vssd1 vssd1 vccd1 vccd1 _2312_/CLK
+ sky130_fd_sc_hd__clkbuf_16
XFILLER_0_38_102 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_38_157 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_30_29 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA_hold980_A _2090_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_34_363 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_219 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_208 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_30_580 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
Xhold4 hold4/A vssd1 vssd1 vccd1 vccd1 hold4/X sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_29_124 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_29_146 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_45_628 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_45_617 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_45_606 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_38_680 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_1823_ _1988_/A vssd1 vssd1 vccd1 vccd1 _1823_/Y sky130_fd_sc_hd__inv_2
X_1754_ _2192_/Q _1756_/B vssd1 vssd1 vccd1 vccd1 _1754_/X sky130_fd_sc_hd__and2_1
XFILLER_0_13_503 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_20_40 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
Xhold404 hold456/X vssd1 vssd1 vccd1 vccd1 hold404/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold426 la_data_in[89] vssd1 vssd1 vccd1 vccd1 hold426/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold415 _1217_/X vssd1 vssd1 vccd1 vccd1 hold415/X sky130_fd_sc_hd__dlymetal6s2s_1
XFILLER_0_40_322 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__1591__A2 _1623_/A2 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xhold448 hold452/X vssd1 vssd1 vccd1 vccd1 hold448/X sky130_fd_sc_hd__buf_1
Xhold459 la_data_in[74] vssd1 vssd1 vccd1 vccd1 hold459/X sky130_fd_sc_hd__dlygate4sd3_1
X_1685_ _2113_/Q _1725_/B vssd1 vssd1 vccd1 vccd1 _1685_/X sky130_fd_sc_hd__and2_2
Xhold437 _1493_/X vssd1 vssd1 vccd1 vccd1 hold437/X sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_40_388 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_742 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_731 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_720 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_786 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_775 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_764 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_753 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_2306_ _2328_/CLK _2306_/D _2045_/Y vssd1 vssd1 vccd1 vccd1 _2306_/Q sky130_fd_sc_hd__dfrtp_1
X_2237_ _2238_/CLK _2237_/D _1977_/Y vssd1 vssd1 vccd1 vccd1 _2237_/Q sky130_fd_sc_hd__dfrtp_1
XTAP_797 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__1361__A _1415_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_24_3 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_2168_ _2168_/CLK _2168_/D _1908_/Y vssd1 vssd1 vccd1 vccd1 _2168_/Q sky130_fd_sc_hd__dfrtp_4
X_2099_ _2182_/CLK _2099_/D _1842_/Y vssd1 vssd1 vccd1 vccd1 _2099_/Q sky130_fd_sc_hd__dfrtp_4
XFILLER_0_48_411 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_1119_ hold648/X _1189_/A2 _1189_/B1 _1118_/X vssd1 vssd1 vccd1 vccd1 _2285_/D sky130_fd_sc_hd__a22o_1
XFILLER_0_48_477 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_48_455 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_29_691 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XANTENNA__1300__S _1318_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_51_609 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__1567__C1 hold406/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_31_377 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xhold960 _1351_/X vssd1 vssd1 vccd1 vccd1 _2194_/D sky130_fd_sc_hd__dlygate4sd3_1
Xhold982 _2099_/Q vssd1 vssd1 vccd1 vccd1 hold982/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold971 _2162_/Q vssd1 vssd1 vccd1 vccd1 hold971/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold993 _2078_/Q vssd1 vssd1 vccd1 vccd1 hold993/X sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA__1098__A1 _2115_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_39_422 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XANTENNA__1210__S _1252_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__1270__A1 _2221_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xoutput509 hold651/X vssd1 vssd1 vccd1 vccd1 la_data_out[94] sky130_fd_sc_hd__buf_12
XFILLER_0_22_333 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_22_344 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_1470_ hold8/X _2151_/Q hold80/X vssd1 vssd1 vccd1 vccd1 hold9/A sky130_fd_sc_hd__mux2_1
X_2022_ _2026_/A vssd1 vssd1 vccd1 vccd1 _2022_/Y sky130_fd_sc_hd__inv_2
XFILLER_0_49_208 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_57_252 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__1261__A1 _2224_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_1806_ _1808_/D _1806_/B _1806_/C _1808_/C vssd1 vssd1 vccd1 vccd1 _1807_/B sky130_fd_sc_hd__or4b_1
XFILLER_0_13_300 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_26_661 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
Xhold201 hold239/X vssd1 vssd1 vccd1 vccd1 hold201/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold212 _1372_/X vssd1 vssd1 vccd1 vccd1 _2187_/D sky130_fd_sc_hd__dlygate4sd3_1
Xhold234 la_data_in[13] vssd1 vssd1 vccd1 vccd1 hold234/X sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_13_366 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
Xhold223 _1361_/X vssd1 vssd1 vccd1 vccd1 hold223/X sky130_fd_sc_hd__dlymetal6s2s_1
X_1737_ _2175_/Q _1766_/B vssd1 vssd1 vccd1 vccd1 _1737_/X sky130_fd_sc_hd__and2_2
XFILLER_0_40_141 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
Xhold245 _1569_/X vssd1 vssd1 vccd1 vccd1 hold245/X sky130_fd_sc_hd__dlygate4sd3_1
X_1668_ _2096_/Q _1677_/B vssd1 vssd1 vccd1 vccd1 _1668_/X sky130_fd_sc_hd__and2_1
Xhold278 la_data_in[30] vssd1 vssd1 vccd1 vccd1 hold278/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold256 la_data_in[28] vssd1 vssd1 vccd1 vccd1 hold256/X sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_13_388 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
Xhold267 _1293_/X vssd1 vssd1 vccd1 vccd1 hold267/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold289 hold289/A vssd1 vssd1 vccd1 vccd1 _1358_/B sky130_fd_sc_hd__dlygate4sd3_1
X_1599_ input71/X _1619_/A2 _1619_/B1 _2087_/Q hold512/X vssd1 vssd1 vccd1 vccd1 _1599_/X
+ sky130_fd_sc_hd__a221o_1
XTAP_561 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_550 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_572 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_583 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_594 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_56_91 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA_fanout564_A _1527_/A2 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__1030__S _1094_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_36_458 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_36_469 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_51_417 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_17_661 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA_clkbuf_leaf_21_wb_clk_i_A clkbuf_1_1__f_wb_clk_i/X vssd1 vssd1 vccd1 vccd1
+ sky130_fd_sc_hd__diode_2
XFILLER_0_16_193 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__1555__A2 _1637_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xhold790 _2150_/Q vssd1 vssd1 vccd1 vccd1 hold790/X sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA__1491__A1 _1491_/A1 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_54_211 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_0970_ _0977_/C _0977_/D hold35/X _0977_/B vssd1 vssd1 vccd1 vccd1 _0970_/X sky130_fd_sc_hd__and4b_1
XFILLER_0_39_274 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_39_285 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_54_233 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_54_222 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_27_458 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_54_277 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
Xoutput306 _1781_/X vssd1 vssd1 vccd1 vccd1 data_out[139] sky130_fd_sc_hd__buf_12
Xoutput317 _1791_/X vssd1 vssd1 vccd1 vccd1 data_out[149] sky130_fd_sc_hd__buf_12
Xoutput339 _1663_/X vssd1 vssd1 vccd1 vccd1 data_out[21] sky130_fd_sc_hd__buf_12
X_1522_ hold392/X _2125_/Q hold80/X vssd1 vssd1 vccd1 vccd1 _1522_/X sky130_fd_sc_hd__mux2_1
Xoutput328 _1801_/X vssd1 vssd1 vccd1 vccd1 data_out[159] sky130_fd_sc_hd__buf_12
X_1453_ _1453_/A _1453_/B _1453_/C _1453_/D vssd1 vssd1 vccd1 vccd1 _1453_/X sky130_fd_sc_hd__or4_1
XANTENNA__1904__A _1913_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_1384_ _1383_/X hold955/X _1435_/S vssd1 vssd1 vccd1 vccd1 _2183_/D sky130_fd_sc_hd__mux2_1
X_2005_ _2034_/A vssd1 vssd1 vccd1 vccd1 _2005_/Y sky130_fd_sc_hd__inv_2
XFILLER_0_9_113 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_45_244 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_42_93 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_18_447 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_5_330 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_14_642 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_41_461 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_5_385 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_14_653 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_14_675 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_41_472 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_13_174 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__1537__A2 _1197_/D vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xfanout533 _1022_/X vssd1 vssd1 vccd1 vccd1 _1097_/A2 sky130_fd_sc_hd__clkbuf_4
Xfanout522 hold26/X vssd1 vssd1 vccd1 vccd1 _1435_/S sky130_fd_sc_hd__buf_6
Xfanout555 _1023_/Y vssd1 vssd1 vccd1 vccd1 _1157_/B1 sky130_fd_sc_hd__clkbuf_4
Xfanout544 _1641_/Y vssd1 vssd1 vccd1 vccd1 _1724_/B sky130_fd_sc_hd__clkbuf_4
Xfanout566 _1527_/A2 vssd1 vssd1 vccd1 vccd1 _1529_/A2 sky130_fd_sc_hd__buf_4
Xfanout599 input262/X vssd1 vssd1 vccd1 vccd1 _1913_/A sky130_fd_sc_hd__clkbuf_8
Xfanout588 _1038_/S vssd1 vssd1 vccd1 vccd1 _1112_/S sky130_fd_sc_hd__buf_4
XTAP_391 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_380 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xfanout577 _1527_/B1 vssd1 vssd1 vccd1 vccd1 _1541_/B1 sky130_fd_sc_hd__buf_4
XANTENNA__1170__A0 _2171_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XPHY_20 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_31 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_42 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__1473__A1 _1473_/A1 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XPHY_53 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_64 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_97 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_86 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_75 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_37_712 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_52_704 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_24_417 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_51_225 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_20_601 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__1724__A _2162_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_47_49 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__1161__B1 _1189_/B1 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_59_369 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_28_701 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XANTENNA_18 la_data_in[51] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_27_222 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_0953_ _0992_/A vssd1 vssd1 vccd1 vccd1 _0953_/Y sky130_fd_sc_hd__inv_2
XFILLER_0_27_266 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_42_225 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_30_409 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__1519__A2 _1519_/A2 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_50_291 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_1505_ _1505_/A1 _1519_/A2 _1519_/B1 _2134_/Q hold475/X vssd1 vssd1 vccd1 vccd1 _1505_/X
+ sky130_fd_sc_hd__a221o_1
XFILLER_0_2_377 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_1436_ _1445_/A _1436_/B vssd1 vssd1 vccd1 vccd1 _1436_/X sky130_fd_sc_hd__and2_1
XANTENNA__1152__A0 _2180_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_1367_ _1415_/A _1367_/B vssd1 vssd1 vccd1 vccd1 _1367_/X sky130_fd_sc_hd__and2_1
XFILLER_0_37_60 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_1298_ _1310_/A _1298_/B vssd1 vssd1 vccd1 vccd1 _1298_/X sky130_fd_sc_hd__and2_1
XFILLER_0_38_509 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_46_542 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_46_531 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_46_520 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA_fanout527_A _1157_/A2 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_18_211 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_18_233 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_21_409 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__1143__B1 _1189_/B1 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__1446__B2 _2163_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__1446__A1 _1446_/A1 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_49_380 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__1719__A _2147_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xinput16 data_in[113] vssd1 vssd1 vccd1 vccd1 input16/X sky130_fd_sc_hd__clkbuf_1
Xinput27 data_in[123] vssd1 vssd1 vccd1 vccd1 input27/X sky130_fd_sc_hd__buf_1
XFILLER_0_3_108 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_37_597 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
Xinput38 data_in[133] vssd1 vssd1 vccd1 vccd1 input38/X sky130_fd_sc_hd__buf_1
Xinput49 data_in[143] vssd1 vssd1 vccd1 vccd1 input49/X sky130_fd_sc_hd__buf_1
XFILLER_0_58_15 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_2270_ _2296_/CLK _2270_/D _2009_/Y vssd1 vssd1 vccd1 vccd1 _2270_/Q sky130_fd_sc_hd__dfrtp_1
X_1221_ input64/X _1503_/A2 _1503_/B1 _2238_/Q hold515/X vssd1 vssd1 vccd1 vccd1 _1221_/X
+ sky130_fd_sc_hd__a221o_1
XANTENNA__1134__A0 _2189_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_1152_ _2180_/Q _2088_/Q _1178_/S vssd1 vssd1 vccd1 vccd1 _1152_/X sky130_fd_sc_hd__mux2_1
X_1083_ _2303_/Q _1095_/A2 _1095_/B1 _1082_/X vssd1 vssd1 vccd1 vccd1 _1083_/X sky130_fd_sc_hd__a22o_1
XANTENNA__1437__B2 _2166_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_28_531 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_1985_ _1988_/A vssd1 vssd1 vccd1 vccd1 _1985_/Y sky130_fd_sc_hd__inv_2
XFILLER_0_16_704 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_28_586 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_15_225 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_31_707 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_43_589 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_2_141 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__1364__A _1415_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_54_3 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_11_497 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_1419_ _1419_/A1 _1198_/A _1545_/B1 _2172_/Q hold101/X vssd1 vssd1 vccd1 vccd1 _1419_/X
+ sky130_fd_sc_hd__a221o_1
XANTENNA__1125__B1 _1183_/B1 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__1303__S _1318_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__1428__B2 _2169_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_38_317 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_19_542 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_53_309 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_34_501 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_46_394 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__1600__A1 _2086_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_34_567 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_34_589 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_28_29 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__1116__A0 _2198_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__1213__S _1252_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__1419__B2 _2172_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_44_309 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_1770_ _2208_/Q _1804_/B vssd1 vssd1 vccd1 vccd1 _1770_/X sky130_fd_sc_hd__and2_1
XFILLER_0_52_331 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_25_545 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
Xhold608 hold736/X vssd1 vssd1 vccd1 vccd1 hold608/X sky130_fd_sc_hd__buf_1
XFILLER_0_52_397 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
Xhold619 _1101_/X vssd1 vssd1 vccd1 vccd1 _2294_/D sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_0_612 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_2322_ _2322_/CLK _2322_/D _2061_/Y vssd1 vssd1 vccd1 vccd1 _2322_/Q sky130_fd_sc_hd__dfrtp_1
XFILLER_0_20_261 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_2253_ _2269_/CLK _2253_/D _1992_/Y vssd1 vssd1 vccd1 vccd1 _2253_/Q sky130_fd_sc_hd__dfrtp_1
XANTENNA__1912__A _1913_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_2184_ _2194_/CLK _2184_/D _1924_/Y vssd1 vssd1 vccd1 vccd1 _2184_/Q sky130_fd_sc_hd__dfrtp_4
X_1204_ hold38/X _1204_/B hold24/X vssd1 vssd1 vccd1 vccd1 hold39/A sky130_fd_sc_hd__or3_1
X_1135_ hold614/X _1157_/A2 _1183_/B1 _1134_/X vssd1 vssd1 vccd1 vccd1 _2277_/D sky130_fd_sc_hd__a22o_1
Xclkbuf_0_wb_clk_i wb_clk_i vssd1 vssd1 vccd1 vccd1 clkbuf_0_wb_clk_i/X sky130_fd_sc_hd__clkbuf_16
X_1066_ _2223_/Q _2131_/Q _1086_/S vssd1 vssd1 vccd1 vccd1 _1066_/X sky130_fd_sc_hd__mux2_1
XFILLER_0_8_701 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_34_83 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_47_169 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_35_309 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_7_266 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_1968_ _1982_/A vssd1 vssd1 vccd1 vccd1 _1968_/Y sky130_fd_sc_hd__inv_2
XFILLER_0_43_364 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_1899_ _1949_/A vssd1 vssd1 vccd1 vccd1 _1899_/Y sky130_fd_sc_hd__inv_2
XFILLER_0_16_589 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA_fanout594_A _0952_/Y vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xinput217 hold468/X vssd1 vssd1 vccd1 vccd1 hold469/A sky130_fd_sc_hd__buf_1
Xinput206 hold139/X vssd1 vssd1 vccd1 vccd1 hold140/A sky130_fd_sc_hd__clkbuf_1
Xinput228 hold357/X vssd1 vssd1 vccd1 vccd1 hold358/A sky130_fd_sc_hd__clkbuf_1
Xinput239 hold229/X vssd1 vssd1 vccd1 vccd1 hold230/A sky130_fd_sc_hd__clkbuf_1
XFILLER_0_39_626 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_39_659 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_53_139 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_53_117 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_47_670 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_34_320 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XANTENNA__1585__B1 _1623_/B1 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_hold973_A _2091_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_209 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__1732__A _2170_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_55_38 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
Xhold5 la_data_in[81] vssd1 vssd1 vccd1 vccd1 hold5/X sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_29_169 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_44_139 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_1822_ _1988_/A vssd1 vssd1 vccd1 vccd1 _1822_/Y sky130_fd_sc_hd__inv_2
XFILLER_0_38_670 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_37_191 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_1753_ _2191_/Q _1756_/B vssd1 vssd1 vccd1 vccd1 _1753_/X sky130_fd_sc_hd__and2_1
XFILLER_0_13_515 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_25_386 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
Xhold405 _1806_/B vssd1 vssd1 vccd1 vccd1 _1349_/B sky130_fd_sc_hd__dlygate4sd3_1
Xhold427 hold427/A vssd1 vssd1 vccd1 vccd1 _1453_/B sky130_fd_sc_hd__buf_1
XFILLER_0_20_85 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_1684_ _2112_/Q _1725_/B vssd1 vssd1 vccd1 vccd1 _1684_/X sky130_fd_sc_hd__and2_1
Xhold416 _1218_/X vssd1 vssd1 vccd1 vccd1 hold416/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold449 hold449/A vssd1 vssd1 vccd1 vccd1 _1277_/B sky130_fd_sc_hd__dlygate4sd3_1
Xhold438 _1494_/X vssd1 vssd1 vccd1 vccd1 _2139_/D sky130_fd_sc_hd__dlygate4sd3_1
XTAP_710 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_21_581 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_743 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_732 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_721 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_29_61 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_776 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_765 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_754 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_2305_ _2328_/CLK _2305_/D _2044_/Y vssd1 vssd1 vccd1 vccd1 _2305_/Q sky130_fd_sc_hd__dfrtp_1
XANTENNA__1642__A _2070_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_2236_ _2238_/CLK _2236_/D _1976_/Y vssd1 vssd1 vccd1 vccd1 _2236_/Q sky130_fd_sc_hd__dfrtp_1
XTAP_787 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_798 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_17_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_2167_ _2168_/CLK _2167_/D _1907_/Y vssd1 vssd1 vccd1 vccd1 _2167_/Q sky130_fd_sc_hd__dfrtp_4
X_2098_ _2168_/CLK _2098_/D _1841_/Y vssd1 vssd1 vccd1 vccd1 _2098_/Q sky130_fd_sc_hd__dfrtp_4
X_1118_ _2197_/Q _2105_/Q _1156_/S vssd1 vssd1 vccd1 vccd1 _1118_/X sky130_fd_sc_hd__mux2_1
X_1049_ hold594/X _1095_/A2 _1095_/B1 _1048_/X vssd1 vssd1 vccd1 vccd1 _2320_/D sky130_fd_sc_hd__a22o_1
XFILLER_0_0_62 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA_clkbuf_leaf_11_wb_clk_i_A clkbuf_1_1__f_wb_clk_i/X vssd1 vssd1 vccd1 vccd1
+ sky130_fd_sc_hd__diode_2
XANTENNA_fanout607_A _2034_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__1567__B1 _1569_/B1 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_31_345 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_12_581 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__1028__S _1094_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xhold972 _2083_/Q vssd1 vssd1 vccd1 vccd1 hold972/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold961 _2201_/Q vssd1 vssd1 vccd1 vccd1 hold961/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold950 _2106_/Q vssd1 vssd1 vccd1 vccd1 hold950/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold994 _2128_/Q vssd1 vssd1 vccd1 vccd1 hold994/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold983 _2074_/Q vssd1 vssd1 vccd1 vccd1 hold983/X sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_39_434 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_26_128 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_35_673 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_41_109 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_50_643 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__1727__A _2165_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_35_695 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_2021_ _2034_/A vssd1 vssd1 vccd1 vccd1 _2021_/Y sky130_fd_sc_hd__inv_2
XANTENNA__1089__A2 _1097_/A2 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_58_710 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_17_128 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_26_640 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_1805_ _1805_/A _1809_/B _1635_/B vssd1 vssd1 vccd1 vccd1 _1806_/C sky130_fd_sc_hd__or3b_1
XFILLER_0_26_673 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_41_632 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xhold202 hold202/A vssd1 vssd1 vccd1 vccd1 _1409_/B sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_13_334 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__1637__A _1637_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_1736_ _2174_/Q _1766_/B vssd1 vssd1 vccd1 vccd1 _1736_/X sky130_fd_sc_hd__and2_1
Xhold224 _1575_/X vssd1 vssd1 vccd1 vccd1 hold224/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold213 hold898/X vssd1 vssd1 vccd1 vccd1 hold213/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold235 hold262/X vssd1 vssd1 vccd1 vccd1 hold263/A sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_13_345 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_1667_ _2095_/Q _1680_/B vssd1 vssd1 vccd1 vccd1 _1667_/X sky130_fd_sc_hd__and2_1
Xhold257 la_data_in[49] vssd1 vssd1 vccd1 vccd1 hold257/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold246 hold251/X vssd1 vssd1 vccd1 vccd1 hold246/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold268 _1294_/X vssd1 vssd1 vccd1 vccd1 _2213_/D sky130_fd_sc_hd__dlygate4sd3_1
X_1598_ _1597_/X hold985/X _1622_/S vssd1 vssd1 vccd1 vccd1 _2087_/D sky130_fd_sc_hd__mux2_1
Xhold279 hold294/X vssd1 vssd1 vccd1 vccd1 hold279/X sky130_fd_sc_hd__dlygate4sd3_1
XTAP_540 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_551 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_562 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_573 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_584 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_595 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_fanout557_A _1097_/B1 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_2219_ _2219_/CLK _2219_/D _1959_/Y vssd1 vssd1 vccd1 vccd1 _2219_/Q sky130_fd_sc_hd__dfrtp_4
XANTENNA__1485__C1 hold422/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_48_253 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_36_415 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_8_350 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_17_673 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_32_643 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xhold780 _1191_/X vssd1 vssd1 vccd1 vccd1 hold780/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold791 _1028_/X vssd1 vssd1 vccd1 vccd1 hold791/X sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_39_297 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_54_267 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_54_256 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xoutput307 _1655_/X vssd1 vssd1 vccd1 vccd1 data_out[13] sky130_fd_sc_hd__buf_12
Xoutput329 _1657_/X vssd1 vssd1 vccd1 vccd1 data_out[15] sky130_fd_sc_hd__buf_12
X_1521_ _1521_/A1 _1527_/A2 _1527_/B1 _2126_/Q hold391/X vssd1 vssd1 vccd1 vccd1 _1521_/X
+ sky130_fd_sc_hd__a221o_1
Xoutput318 _1656_/X vssd1 vssd1 vccd1 vccd1 data_out[14] sky130_fd_sc_hd__buf_12
XFILLER_0_10_315 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_10_348 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_1452_ hold90/X _2159_/Q _1461_/S vssd1 vssd1 vccd1 vccd1 _1452_/X sky130_fd_sc_hd__mux2_1
X_1383_ input5/X _1533_/A2 _1533_/B1 _2184_/Q hold529/X vssd1 vssd1 vccd1 vccd1 _1383_/X
+ sky130_fd_sc_hd__a221o_1
XANTENNA__1920__A _1922_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_2004_ _2008_/A vssd1 vssd1 vccd1 vccd1 _2004_/Y sky130_fd_sc_hd__inv_2
XFILLER_0_42_61 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_42_50 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_45_223 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_9_169 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_45_278 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_45_289 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__1367__A _1415_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_14_610 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_26_481 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_1719_ _2147_/Q _1756_/B vssd1 vssd1 vccd1 vccd1 _1719_/X sky130_fd_sc_hd__and2_1
Xfanout523 hold26/X vssd1 vssd1 vccd1 vccd1 _1372_/S sky130_fd_sc_hd__clkbuf_4
Xfanout556 _1097_/B1 vssd1 vssd1 vccd1 vccd1 _1095_/B1 sky130_fd_sc_hd__buf_4
Xfanout534 hold80/X vssd1 vssd1 vccd1 vccd1 _1632_/S sky130_fd_sc_hd__clkbuf_8
Xfanout545 _1766_/B vssd1 vssd1 vccd1 vccd1 _1804_/B sky130_fd_sc_hd__clkbuf_4
XANTENNA__1306__S _1318_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xfanout567 _1003_/Y vssd1 vssd1 vccd1 vccd1 _1527_/A2 sky130_fd_sc_hd__buf_4
XTAP_370 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_392 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_381 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__1170__A1 _2079_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xfanout578 _1529_/B1 vssd1 vssd1 vccd1 vccd1 _1533_/B1 sky130_fd_sc_hd__buf_4
Xfanout589 _1094_/S vssd1 vssd1 vccd1 vccd1 _1086_/S sky130_fd_sc_hd__clkbuf_8
XPHY_21 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_10 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_32 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_43 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_54 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_65 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_98 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_87 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_76 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_51_248 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XANTENNA__1724__B _1724_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__1216__S _1252_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__1740__A _2178_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_59_337 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_28_713 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA_19 hold275/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_0952_ _2249_/Q vssd1 vssd1 vccd1 vccd1 _0952_/Y sky130_fd_sc_hd__inv_2
XFILLER_0_43_705 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_27_278 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_2_334 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_23_484 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_2_389 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_1504_ _1503_/X _2134_/Q _1504_/S vssd1 vssd1 vccd1 vccd1 _1504_/X sky130_fd_sc_hd__mux2_1
X_1435_ hold282/X hold979/X _1435_/S vssd1 vssd1 vccd1 vccd1 _2166_/D sky130_fd_sc_hd__mux2_1
XANTENNA__1152__A1 _2088_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_1366_ _1365_/X hold926/X _1372_/S vssd1 vssd1 vccd1 vccd1 _2189_/D sky130_fd_sc_hd__mux2_1
XANTENNA__1650__A _2078_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_1297_ hold165/X _2212_/Q _1318_/S vssd1 vssd1 vccd1 vccd1 _1297_/X sky130_fd_sc_hd__mux2_1
XFILLER_0_19_713 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_18_245 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_34_705 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_14_451 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_41_281 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xclkbuf_leaf_15_wb_clk_i clkbuf_1_1__f_wb_clk_i/X vssd1 vssd1 vccd1 vccd1 _2300_/CLK
+ sky130_fd_sc_hd__clkbuf_16
XFILLER_0_56_307 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xinput28 data_in[124] vssd1 vssd1 vccd1 vccd1 input28/X sky130_fd_sc_hd__buf_1
Xinput17 data_in[114] vssd1 vssd1 vccd1 vccd1 input17/X sky130_fd_sc_hd__clkbuf_1
Xinput39 data_in[134] vssd1 vssd1 vccd1 vccd1 input39/X sky130_fd_sc_hd__buf_1
XFILLER_0_20_421 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XANTENNA__1735__A _2173_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_32_292 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_1220_ _1277_/A _1220_/B vssd1 vssd1 vccd1 vccd1 _1220_/X sky130_fd_sc_hd__and2_1
XANTENNA__1134__A1 _2097_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_1151_ hold626/X _1183_/A2 _1183_/B1 _1150_/X vssd1 vssd1 vccd1 vccd1 _2269_/D sky130_fd_sc_hd__a22o_1
X_1082_ _2215_/Q _2123_/Q _1086_/S vssd1 vssd1 vccd1 vccd1 _1082_/X sky130_fd_sc_hd__mux2_1
X_1984_ _1988_/A vssd1 vssd1 vccd1 vccd1 _1984_/Y sky130_fd_sc_hd__inv_2
XFILLER_0_43_535 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_15_215 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__1070__A0 _2221_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_15_237 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_15_259 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_43_579 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_11_410 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_23_292 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__1645__A _2073_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_2_197 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_47_3 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_1418_ _1445_/A _1418_/B vssd1 vssd1 vccd1 vccd1 _1418_/X sky130_fd_sc_hd__and2_1
X_1349_ _1349_/A _1349_/B vssd1 vssd1 vccd1 vccd1 _1349_/X sky130_fd_sc_hd__and2_1
XANTENNA__1428__A2 _1569_/A2 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_38_307 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_19_554 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__1061__B1 _1095_/B1 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_21_229 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xoutput490 hold593/X vssd1 vssd1 vccd1 vccd1 la_data_out[75] sky130_fd_sc_hd__buf_12
XANTENNA__1116__A1 _2106_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_25_502 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_25_557 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_52_365 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
Xhold609 _1161_/X vssd1 vssd1 vccd1 vccd1 _2264_/D sky130_fd_sc_hd__dlygate4sd3_1
X_2321_ _2330_/CLK _2321_/D _2060_/Y vssd1 vssd1 vccd1 vccd1 _2321_/Q sky130_fd_sc_hd__dfrtp_1
X_2252_ _2291_/CLK _2252_/D _1991_/Y vssd1 vssd1 vccd1 vccd1 _2252_/Q sky130_fd_sc_hd__dfrtp_1
X_1203_ _0986_/Y _1192_/B hold23/X _1202_/Y vssd1 vssd1 vccd1 vccd1 hold24/A sky130_fd_sc_hd__a31o_1
X_2183_ _2194_/CLK _2183_/D _1923_/Y vssd1 vssd1 vccd1 vccd1 _2183_/Q sky130_fd_sc_hd__dfrtp_4
X_1134_ _2189_/Q _2097_/Q _1156_/S vssd1 vssd1 vccd1 vccd1 _1134_/X sky130_fd_sc_hd__mux2_1
XFILLER_0_18_96 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_1065_ hold651/X _1095_/A2 _1095_/B1 _1064_/X vssd1 vssd1 vccd1 vccd1 _2312_/D sky130_fd_sc_hd__a22o_1
XFILLER_0_19_7 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_34_62 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_8_713 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_7_223 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_7_201 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_28_351 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_7_256 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_50_83 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_43_343 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_16_568 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_1967_ _1979_/A vssd1 vssd1 vccd1 vccd1 _1967_/Y sky130_fd_sc_hd__inv_2
XFILLER_0_43_387 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_1898_ _1949_/A vssd1 vssd1 vccd1 vccd1 _1898_/Y sky130_fd_sc_hd__inv_2
XANTENNA_fanout587_A _1112_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xinput207 hold145/X vssd1 vssd1 vccd1 vccd1 hold146/A sky130_fd_sc_hd__buf_1
Xinput218 hold461/X vssd1 vssd1 vccd1 vccd1 hold462/A sky130_fd_sc_hd__clkbuf_1
Xinput229 hold434/X vssd1 vssd1 vccd1 vccd1 hold435/A sky130_fd_sc_hd__clkbuf_1
XFILLER_0_38_137 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_39_638 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_19_384 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_34_332 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_22_527 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__1585__B2 _2094_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_22_549 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_34_387 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA_hold966_A _2181_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_30_560 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xhold6 hold6/A vssd1 vssd1 vccd1 vccd1 hold6/X sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_57_446 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_1821_ _1852_/A vssd1 vssd1 vccd1 vccd1 _1821_/Y sky130_fd_sc_hd__inv_2
XFILLER_0_53_685 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_52_162 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_1752_ _2190_/Q _1761_/B vssd1 vssd1 vccd1 vccd1 _1752_/X sky130_fd_sc_hd__and2_1
XFILLER_0_52_195 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_52_173 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
Xhold417 _1219_/X vssd1 vssd1 vccd1 vccd1 _2238_/D sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_20_53 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_1683_ _2111_/Q _1725_/B vssd1 vssd1 vccd1 vccd1 _1683_/X sky130_fd_sc_hd__and2_2
Xhold406 _1349_/X vssd1 vssd1 vccd1 vccd1 hold406/X sky130_fd_sc_hd__dlymetal6s2s_1
Xhold428 _0980_/X vssd1 vssd1 vccd1 vccd1 hold428/X sky130_fd_sc_hd__clkdlybuf4s25_1
Xhold439 la_data_in[54] vssd1 vssd1 vccd1 vccd1 hold439/X sky130_fd_sc_hd__dlygate4sd3_1
XTAP_700 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__1923__A _1941_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_733 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_711 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_722 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_777 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_766 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_755 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_744 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_2304_ _2328_/CLK _2304_/D _2043_/Y vssd1 vssd1 vccd1 vccd1 _2304_/Q sky130_fd_sc_hd__dfrtp_1
XTAP_788 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_799 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_2235_ _2238_/CLK _2235_/D _1975_/Y vssd1 vssd1 vccd1 vccd1 _2235_/Q sky130_fd_sc_hd__dfrtp_1
XANTENNA__1642__B _1725_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_2166_ _2177_/CLK _2166_/D _1906_/Y vssd1 vssd1 vccd1 vccd1 _2166_/Q sky130_fd_sc_hd__dfrtp_4
X_1117_ hold649/X _1183_/A2 _1183_/B1 _1116_/X vssd1 vssd1 vccd1 vccd1 _2286_/D sky130_fd_sc_hd__a22o_1
X_2097_ _2168_/CLK _2097_/D _1840_/Y vssd1 vssd1 vccd1 vccd1 _2097_/Q sky130_fd_sc_hd__dfrtp_4
XFILLER_0_45_94 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_1048_ _2232_/Q _2140_/Q _1094_/S vssd1 vssd1 vccd1 vccd1 _1048_/X sky130_fd_sc_hd__mux2_1
XFILLER_0_48_446 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_35_118 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_44_641 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_16_332 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_16_365 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_16_376 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XANTENNA__1567__B2 _2103_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_clkbuf_leaf_7_wb_clk_i_A clkbuf_leaf_9_wb_clk_i/A vssd1 vssd1 vccd1 vccd1
+ sky130_fd_sc_hd__diode_2
Xhold940 _2104_/Q vssd1 vssd1 vccd1 vccd1 hold940/X sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA__1309__S _1318_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_31_357 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
Xhold973 _2091_/Q vssd1 vssd1 vccd1 vccd1 hold973/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold962 _2098_/Q vssd1 vssd1 vccd1 vccd1 hold962/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold951 _2074_/Q vssd1 vssd1 vccd1 vccd1 hold951/X sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA__1833__A _1922_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xhold984 _2165_/Q vssd1 vssd1 vccd1 vccd1 hold984/X sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_39_402 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_39_446 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_39_468 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_35_685 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__1558__A1 _2107_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_34_162 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_34_195 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__1219__S _1252_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_50_699 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__1743__A _2181_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_2020_ _2033_/A vssd1 vssd1 vccd1 vccd1 _2020_/Y sky130_fd_sc_hd__inv_2
XFILLER_0_15_20 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_15_64 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_57_243 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_45_405 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_45_449 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XANTENNA__1918__A _1941_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_31_52 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_1804_ _2242_/Q _1804_/B vssd1 vssd1 vccd1 vccd1 _1804_/X sky130_fd_sc_hd__and2_1
XANTENNA__1637__B _1637_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__1549__B2 _2112_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_26_685 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_1735_ _2173_/Q _1766_/B vssd1 vssd1 vccd1 vccd1 _1735_/X sky130_fd_sc_hd__and2_1
XFILLER_0_41_655 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xhold225 hold302/X vssd1 vssd1 vccd1 vccd1 hold225/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold214 la_data_in[79] vssd1 vssd1 vccd1 vccd1 hold214/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold203 _1409_/X vssd1 vssd1 vccd1 vccd1 hold203/X sky130_fd_sc_hd__buf_1
XFILLER_0_40_154 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
Xhold236 hold236/A vssd1 vssd1 vccd1 vccd1 _1364_/B sky130_fd_sc_hd__dlygate4sd3_1
Xhold247 hold247/A vssd1 vssd1 vccd1 vccd1 _1367_/B sky130_fd_sc_hd__dlygate4sd3_1
Xhold269 hold424/X vssd1 vssd1 vccd1 vccd1 hold269/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold258 _1300_/X vssd1 vssd1 vccd1 vccd1 _2211_/D sky130_fd_sc_hd__dlygate4sd3_1
X_1666_ _2094_/Q _1680_/B vssd1 vssd1 vccd1 vccd1 _1666_/X sky130_fd_sc_hd__and2_1
X_1597_ input72/X _1619_/A2 _1619_/B1 _2088_/Q _1394_/X vssd1 vssd1 vccd1 vccd1 _1597_/X
+ sky130_fd_sc_hd__a221o_1
XANTENNA__1653__A _2081_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_530 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_541 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_552 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_563 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_574 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_585 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_596 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_2218_ _2223_/CLK _2218_/D _1958_/Y vssd1 vssd1 vccd1 vccd1 _2218_/Q sky130_fd_sc_hd__dfrtp_4
X_2149_ _2322_/CLK _2149_/D _1892_/Y vssd1 vssd1 vccd1 vccd1 _2149_/Q sky130_fd_sc_hd__dfrtp_1
XANTENNA__1485__B1 _1503_/B1 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_8_362 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_51_408 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_8_384 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_17_685 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_32_611 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_32_622 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_31_165 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xhold770 hold770/A vssd1 vssd1 vccd1 vccd1 hold770/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold781 la_data_in[90] vssd1 vssd1 vccd1 vccd1 hold781/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold792 _2116_/Q vssd1 vssd1 vccd1 vccd1 hold792/X sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA_hold929_A _2100_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_59_508 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__1502__S _1504_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__1738__A _2176_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xoutput308 _1782_/X vssd1 vssd1 vccd1 vccd1 data_out[140] sky130_fd_sc_hd__buf_12
XFILLER_0_23_644 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_1520_ _1519_/X _2126_/Q _1520_/S vssd1 vssd1 vccd1 vccd1 _1520_/X sky130_fd_sc_hd__mux2_1
Xoutput319 _1792_/X vssd1 vssd1 vccd1 vccd1 data_out[150] sky130_fd_sc_hd__buf_12
XFILLER_0_10_305 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_22_165 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_50_496 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_1451_ _0974_/X _1192_/B hold89/X vssd1 vssd1 vccd1 vccd1 _1451_/X sky130_fd_sc_hd__a21o_1
X_1382_ _1394_/A _1382_/B vssd1 vssd1 vccd1 vccd1 _1382_/X sky130_fd_sc_hd__and2_1
XFILLER_0_26_41 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_2003_ _2008_/A vssd1 vssd1 vccd1 vccd1 _2003_/Y sky130_fd_sc_hd__inv_2
XFILLER_0_26_74 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_26_85 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_58_530 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__1648__A _2076_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_14_622 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_14_666 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_1718_ _2146_/Q _1761_/B vssd1 vssd1 vccd1 vccd1 _1718_/X sky130_fd_sc_hd__and2_1
XFILLER_0_14_699 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_1649_ _2077_/Q _1677_/B vssd1 vssd1 vccd1 vccd1 _1649_/X sky130_fd_sc_hd__and2_1
Xfanout524 hold26/X vssd1 vssd1 vccd1 vccd1 _1318_/S sky130_fd_sc_hd__clkbuf_8
Xfanout557 _1097_/B1 vssd1 vssd1 vccd1 vccd1 _1057_/B1 sky130_fd_sc_hd__clkbuf_4
XTAP_360 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xfanout546 _1792_/B vssd1 vssd1 vccd1 vccd1 _1766_/B sky130_fd_sc_hd__clkbuf_4
Xfanout535 hold81/X vssd1 vssd1 vccd1 vccd1 _1622_/S sky130_fd_sc_hd__clkbuf_8
XTAP_382 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_371 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_393 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xfanout579 _1527_/B1 vssd1 vssd1 vccd1 vccd1 _1529_/B1 sky130_fd_sc_hd__clkbuf_8
Xfanout568 _1463_/B vssd1 vssd1 vccd1 vccd1 _1503_/A2 sky130_fd_sc_hd__clkbuf_8
XPHY_22 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_11 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_33 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_44 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_55 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_88 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_66 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_77 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_99 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_36_224 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_24_408 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_44_290 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_32_441 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__1161__A2 _1189_/A2 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__1740__B _1761_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__1621__B1 _1623_/B1 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_23_474 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_1503_ _1503_/A1 _1503_/A2 _1503_/B1 _2135_/Q hold317/X vssd1 vssd1 vccd1 vccd1 _1503_/X
+ sky130_fd_sc_hd__a221o_1
X_1434_ _1434_/A1 _1569_/A2 _1569_/B1 _2167_/Q hold281/X vssd1 vssd1 vccd1 vccd1 _1434_/X
+ sky130_fd_sc_hd__a221o_1
XANTENNA__1931__A _1957_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_1365_ input11/X _1529_/A2 _1533_/B1 _2190_/Q hold237/X vssd1 vssd1 vccd1 vccd1 _1365_/X
+ sky130_fd_sc_hd__a221o_1
XFILLER_0_37_51 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_1296_ input37/X _1529_/A2 _1529_/B1 _2213_/Q hold164/X vssd1 vssd1 vccd1 vccd1 _1296_/X
+ sky130_fd_sc_hd__a221o_1
XFILLER_0_46_533 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_46_555 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_5_140 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_14_485 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__2002__A _2002_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__1841__A _1922_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_190 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__1143__A2 _1189_/A2 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__1052__S _1094_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_49_360 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_25_706 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
Xinput18 data_in[115] vssd1 vssd1 vccd1 vccd1 input18/X sky130_fd_sc_hd__clkbuf_1
XFILLER_0_52_525 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__1603__B1 _1623_/B1 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xinput29 data_in[125] vssd1 vssd1 vccd1 vccd1 input29/X sky130_fd_sc_hd__buf_1
XFILLER_0_24_249 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_20_433 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_20_477 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_1150_ _2181_/Q _2089_/Q _1178_/S vssd1 vssd1 vccd1 vccd1 _1150_/X sky130_fd_sc_hd__mux2_1
XANTENNA__1751__A _2189_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_59_113 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_1081_ _2304_/Q _1095_/A2 _1095_/B1 _1080_/X vssd1 vssd1 vccd1 vccd1 _1081_/X sky130_fd_sc_hd__a22o_1
XFILLER_0_28_533 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_1983_ _1988_/A vssd1 vssd1 vccd1 vccd1 _1983_/Y sky130_fd_sc_hd__inv_2
XFILLER_0_55_385 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_43_503 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_43_569 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_43_547 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_15_249 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_11_400 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__1926__A _1941_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_11_422 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_2_165 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_23_260 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__1645__B _1725_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_48_83 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_1417_ _1416_/X _2172_/Q hold27/X vssd1 vssd1 vccd1 vccd1 _1417_/X sky130_fd_sc_hd__mux2_1
XANTENNA__1661__A _2089_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__1125__A2 _1183_/A2 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_1348_ hold107/X hold978/X _1372_/S vssd1 vssd1 vccd1 vccd1 _2195_/D sky130_fd_sc_hd__mux2_1
X_1279_ hold451/X hold957/X _1318_/S vssd1 vssd1 vccd1 vccd1 _2218_/D sky130_fd_sc_hd__mux2_1
XANTENNA_fanout532_A _1097_/A2 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_19_500 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_19_522 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_19_599 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__1597__C1 _1394_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_22_709 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_34_547 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_6_493 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_21_219 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
Xoutput480 hold647/X vssd1 vssd1 vccd1 vccd1 la_data_out[65] sky130_fd_sc_hd__buf_12
Xoutput491 hold618/X vssd1 vssd1 vccd1 vccd1 la_data_out[76] sky130_fd_sc_hd__buf_12
XFILLER_0_29_308 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__1510__S _1520_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_25_525 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_4_419 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_37_396 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__1746__A _2184_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_52_377 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XANTENNA_output451_A hold628/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_2320_ _2328_/CLK _2320_/D _2059_/Y vssd1 vssd1 vccd1 vccd1 _2320_/Q sky130_fd_sc_hd__dfrtp_1
X_2251_ _2251_/CLK _2251_/D _1990_/Y vssd1 vssd1 vccd1 vccd1 _2251_/Q sky130_fd_sc_hd__dfrtp_1
X_1202_ _2248_/Q _1202_/A2 _1193_/Y vssd1 vssd1 vccd1 vccd1 _1202_/Y sky130_fd_sc_hd__a21oi_1
XFILLER_0_18_53 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_2182_ _2182_/CLK _2182_/D _1922_/Y vssd1 vssd1 vccd1 vccd1 _2182_/Q sky130_fd_sc_hd__dfrtp_4
X_1133_ _2278_/Q _1183_/A2 _1157_/B1 _1132_/X vssd1 vssd1 vccd1 vccd1 _1133_/X sky130_fd_sc_hd__a22o_1
X_1064_ _2224_/Q _2132_/Q _1086_/S vssd1 vssd1 vccd1 vccd1 _1064_/X sky130_fd_sc_hd__mux2_1
XANTENNA__1420__S hold27/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xclkbuf_leaf_0_wb_clk_i clkbuf_leaf_9_wb_clk_i/A vssd1 vssd1 vccd1 vccd1 _2173_/CLK
+ sky130_fd_sc_hd__clkbuf_16
XFILLER_0_34_74 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_34_85 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__1291__A1 _2214_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_28_363 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_1966_ _2039_/A vssd1 vssd1 vccd1 vccd1 _1966_/Y sky130_fd_sc_hd__inv_2
XANTENNA__1579__C1 hold248/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_1897_ _2065_/A vssd1 vssd1 vccd1 vccd1 _1897_/Y sky130_fd_sc_hd__inv_2
XFILLER_0_3_430 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__1656__A _2084_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xinput208 hold279/X vssd1 vssd1 vccd1 vccd1 hold280/A sky130_fd_sc_hd__clkbuf_1
Xinput219 hold66/X vssd1 vssd1 vccd1 vccd1 hold67/A sky130_fd_sc_hd__buf_1
XANTENNA__1330__S hold27/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_38_105 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_38_127 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__1282__A1 _2217_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_53_108 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_19_363 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_34_344 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XANTENNA__1034__A1 _2147_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__1585__A2 _1623_/A2 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_22_539 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_34_399 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_30_550 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_30_572 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA_hold959_A _2194_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xhold7 hold7/A vssd1 vssd1 vccd1 vccd1 hold7/X sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA__1240__S _1252_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_45_609 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__1273__A1 _2220_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_1820_ _1852_/A vssd1 vssd1 vccd1 vccd1 _1820_/Y sky130_fd_sc_hd__inv_2
XFILLER_0_38_661 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_38_683 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_25_333 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_52_141 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_1751_ _2189_/Q _1792_/B vssd1 vssd1 vccd1 vccd1 _1751_/X sky130_fd_sc_hd__and2_1
XFILLER_0_25_377 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xhold407 _1567_/X vssd1 vssd1 vccd1 vccd1 hold407/X sky130_fd_sc_hd__dlygate4sd3_1
X_1682_ _2110_/Q _1715_/B vssd1 vssd1 vccd1 vccd1 _1682_/X sky130_fd_sc_hd__and2_1
Xhold418 la_data_in[70] vssd1 vssd1 vccd1 vccd1 hold418/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold429 _0985_/Y vssd1 vssd1 vccd1 vccd1 _0986_/B sky130_fd_sc_hd__dlygate4sd3_1
XTAP_701 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_734 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_712 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_723 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_2303_ _2312_/CLK _2303_/D _2042_/Y vssd1 vssd1 vccd1 vccd1 _2303_/Q sky130_fd_sc_hd__dfrtp_1
XFILLER_0_29_41 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_767 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_756 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_745 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_789 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_778 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_2234_ _2238_/CLK _2234_/D _1974_/Y vssd1 vssd1 vccd1 vccd1 _2234_/Q sky130_fd_sc_hd__dfrtp_1
X_2165_ _2173_/CLK _2165_/D _1905_/Y vssd1 vssd1 vccd1 vccd1 _2165_/Q sky130_fd_sc_hd__dfrtp_4
X_1116_ _2198_/Q _2106_/Q _1178_/S vssd1 vssd1 vccd1 vccd1 _1116_/X sky130_fd_sc_hd__mux2_1
X_2096_ _2168_/CLK _2096_/D _1839_/Y vssd1 vssd1 vccd1 vccd1 _2096_/Q sky130_fd_sc_hd__dfrtp_4
X_1047_ hold595/X _1057_/A2 _1057_/B1 _1046_/X vssd1 vssd1 vccd1 vccd1 _2321_/D sky130_fd_sc_hd__a22o_1
XFILLER_0_28_193 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__1567__A2 _1569_/A2 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_16_344 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_1949_ _1949_/A vssd1 vssd1 vccd1 vccd1 _1949_/Y sky130_fd_sc_hd__inv_2
XFILLER_0_16_388 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
Xhold930 _2119_/Q vssd1 vssd1 vccd1 vccd1 hold930/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold941 _2193_/Q vssd1 vssd1 vccd1 vccd1 hold941/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold963 _2088_/Q vssd1 vssd1 vccd1 vccd1 hold963/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold952 _1624_/X vssd1 vssd1 vccd1 vccd1 _2074_/D sky130_fd_sc_hd__dlygate4sd3_1
Xhold985 _2087_/Q vssd1 vssd1 vccd1 vccd1 hold985/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold974 _2219_/Q vssd1 vssd1 vccd1 vccd1 hold974/X sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_19_160 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_35_631 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_34_141 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_22_347 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_57_222 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_1803_ _2241_/Q _1804_/B vssd1 vssd1 vccd1 vccd1 _1803_/X sky130_fd_sc_hd__and2_1
XANTENNA__1549__A2 _1637_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_25_163 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_1734_ _2172_/Q _1766_/B vssd1 vssd1 vccd1 vccd1 _1734_/X sky130_fd_sc_hd__and2_1
XFILLER_0_26_697 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_40_111 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xhold226 hold226/A vssd1 vssd1 vccd1 vccd1 _1331_/B sky130_fd_sc_hd__dlygate4sd3_1
Xhold215 _1210_/X vssd1 vssd1 vccd1 vccd1 _2241_/D sky130_fd_sc_hd__dlygate4sd3_1
Xhold204 _1607_/X vssd1 vssd1 vccd1 vccd1 hold204/X sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_40_133 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_1665_ _2093_/Q _1680_/B vssd1 vssd1 vccd1 vccd1 _1665_/X sky130_fd_sc_hd__and2_1
Xhold259 hold857/X vssd1 vssd1 vccd1 vccd1 hold259/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold237 _1364_/X vssd1 vssd1 vccd1 vccd1 hold237/X sky130_fd_sc_hd__dlymetal6s2s_1
Xhold248 _1367_/X vssd1 vssd1 vccd1 vccd1 hold248/X sky130_fd_sc_hd__dlymetal6s2s_1
XFILLER_0_40_166 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_1596_ _1595_/X hold963/X _1622_/S vssd1 vssd1 vccd1 vccd1 _2088_/D sky130_fd_sc_hd__mux2_1
XANTENNA__1653__B _1725_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_520 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_531 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_542 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_564 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_553 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_575 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_2217_ _2217_/CLK _2217_/D _1957_/Y vssd1 vssd1 vccd1 vccd1 _2217_/Q sky130_fd_sc_hd__dfrtp_4
XTAP_586 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_597 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_56_94 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_22_3 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XANTENNA__1485__A1 _1485_/A1 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_2148_ _2322_/CLK _2148_/D _1891_/Y vssd1 vssd1 vccd1 vccd1 _2148_/Q sky130_fd_sc_hd__dfrtp_1
X_2079_ _2164_/CLK _2079_/D _1822_/Y vssd1 vssd1 vccd1 vccd1 _2079_/Q sky130_fd_sc_hd__dfrtp_4
XFILLER_0_48_222 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_48_288 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_17_697 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XANTENNA__2005__A _2034_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_32_645 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
Xhold782 _1014_/D vssd1 vssd1 vccd1 vccd1 _0990_/D sky130_fd_sc_hd__dlygate4sd3_1
Xhold771 _2159_/Q vssd1 vssd1 vccd1 vccd1 hold771/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold760 _1196_/X vssd1 vssd1 vccd1 vccd1 hold760/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold793 _2108_/Q vssd1 vssd1 vccd1 vccd1 hold793/X sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA__1173__B1 _1183_/B1 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_52_19 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_54_236 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_54_225 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__1738__B _1761_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_22_133 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
Xoutput309 _1783_/X vssd1 vssd1 vccd1 vccd1 data_out[141] sky130_fd_sc_hd__buf_12
XANTENNA__1754__A _2192_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_1450_ hold2/X hold88/X _1198_/X _1545_/B1 vssd1 vssd1 vccd1 vccd1 hold89/A sky130_fd_sc_hd__a31o_1
X_1381_ _1380_/X hold925/X _1435_/S vssd1 vssd1 vccd1 vccd1 _2184_/D sky130_fd_sc_hd__mux2_1
XANTENNA__1164__A0 _2174_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_2002_ _2002_/A vssd1 vssd1 vccd1 vccd1 _2002_/Y sky130_fd_sc_hd__inv_2
XFILLER_0_58_586 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__1929__A _1941_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_45_203 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_45_225 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_42_74 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_45_247 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_26_472 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__1664__A _2092_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_1717_ _2145_/Q _1798_/B vssd1 vssd1 vccd1 vccd1 _1717_/X sky130_fd_sc_hd__and2_1
XFILLER_0_41_475 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_14_678 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_1648_ _2076_/Q _1677_/B vssd1 vssd1 vccd1 vccd1 _1648_/X sky130_fd_sc_hd__and2_1
Xfanout547 _1761_/B vssd1 vssd1 vccd1 vccd1 _1756_/B sky130_fd_sc_hd__clkbuf_4
X_1579_ input82/X _1619_/A2 _1619_/B1 _2097_/Q hold248/X vssd1 vssd1 vccd1 vccd1 _1579_/X
+ sky130_fd_sc_hd__a221o_1
XANTENNA__1155__B1 _1189_/B1 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_6_96 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_350 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xfanout525 hold26/X vssd1 vssd1 vccd1 vccd1 _1252_/S sky130_fd_sc_hd__buf_6
Xfanout536 hold80/X vssd1 vssd1 vccd1 vccd1 hold81/A sky130_fd_sc_hd__clkbuf_1
Xfanout558 _1023_/Y vssd1 vssd1 vccd1 vccd1 _1097_/B1 sky130_fd_sc_hd__clkbuf_4
XTAP_361 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_383 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_372 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_394 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xfanout569 _1463_/B vssd1 vssd1 vccd1 vccd1 _1495_/A2 sky130_fd_sc_hd__buf_2
XANTENNA_fanout562_A _1569_/A2 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XPHY_12 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_23 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_34 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_45 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_56 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_89 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__1839__A _1922_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XPHY_67 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_78 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__1630__A1 _2071_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_36_247 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_51_206 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_17_483 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_32_464 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_32_497 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__1146__A0 _2183_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xhold590 hold727/X vssd1 vssd1 vccd1 vccd1 hold590/X sky130_fd_sc_hd__clkbuf_2
XANTENNA_hold941_A _2193_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__1749__A _2187_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_12_11 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__1621__B2 _2076_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_12_55 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_2_347 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_1502_ _1501_/X _2135_/Q _1504_/S vssd1 vssd1 vccd1 vccd1 _1502_/X sky130_fd_sc_hd__mux2_1
X_1433_ _1445_/A _1433_/B vssd1 vssd1 vccd1 vccd1 _1433_/X sky130_fd_sc_hd__and2_1
X_1364_ _1415_/A _1364_/B vssd1 vssd1 vccd1 vccd1 _1364_/X sky130_fd_sc_hd__and2_1
X_1295_ _1310_/A _1295_/B vssd1 vssd1 vccd1 vccd1 _1295_/X sky130_fd_sc_hd__and2_1
XANTENNA__1423__S hold27/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_clkbuf_leaf_20_wb_clk_i_A clkbuf_1_1__f_wb_clk_i/X vssd1 vssd1 vccd1 vccd1
+ sky130_fd_sc_hd__diode_2
XFILLER_0_53_73 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__1659__A _2087_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_46_567 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_18_236 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__1612__A1 _2080_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_33_206 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_33_239 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_14_475 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__1128__A0 _2192_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_191 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_180 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__1333__S hold27/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xclkbuf_leaf_24_wb_clk_i clkbuf_leaf_9_wb_clk_i/A vssd1 vssd1 vccd1 vccd1 _2251_/CLK
+ sky130_fd_sc_hd__clkbuf_16
Xinput19 data_in[116] vssd1 vssd1 vccd1 vccd1 input19/X sky130_fd_sc_hd__clkbuf_1
XANTENNA__1603__B2 _2085_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_hold989_A _2111_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_58_29 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__1508__S _1520_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__1119__B1 _1189_/B1 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_20_489 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__1751__B _1792_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__1243__S _1252_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_1080_ _2216_/Q _2124_/Q _1086_/S vssd1 vssd1 vccd1 vccd1 _1080_/X sky130_fd_sc_hd__mux2_1
XFILLER_0_16_707 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_1982_ _1982_/A vssd1 vssd1 vccd1 vccd1 _1982_/Y sky130_fd_sc_hd__inv_2
XFILLER_0_43_526 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_28_589 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_43_559 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_48_51 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_48_40 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__1942__A _1949_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_1416_ _1416_/A1 _1637_/B _1545_/B1 _2173_/Q hold54/X vssd1 vssd1 vccd1 vccd1 _1416_/X
+ sky130_fd_sc_hd__a221o_1
X_1347_ input18/X _1533_/A2 _1533_/B1 _2196_/Q hold106/X vssd1 vssd1 vccd1 vccd1 _1347_/X
+ sky130_fd_sc_hd__a221o_1
XFILLER_0_3_31 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_1278_ input43/X _1519_/A2 _1519_/B1 _2219_/Q hold450/X vssd1 vssd1 vccd1 vccd1 _1278_/X
+ sky130_fd_sc_hd__a221o_1
XFILLER_0_3_86 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_38_309 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_59_670 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_19_545 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA_fanout525_A hold26/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_19_589 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_46_397 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__1061__A2 _1095_/A2 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_42_581 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xoutput470 hold616/X vssd1 vssd1 vccd1 vccd1 la_data_out[55] sky130_fd_sc_hd__buf_12
Xoutput492 hold566/X vssd1 vssd1 vccd1 vccd1 la_data_out[77] sky130_fd_sc_hd__buf_12
Xoutput481 hold643/X vssd1 vssd1 vccd1 vccd1 la_data_out[66] sky130_fd_sc_hd__buf_12
XANTENNA__1521__B1 _1527_/B1 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_37_331 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_52_301 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_52_389 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_33_581 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_0_615 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_20_231 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_20_264 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_2250_ _2291_/CLK _2250_/D _1989_/Y vssd1 vssd1 vccd1 vccd1 _2250_/Q sky130_fd_sc_hd__dfrtp_1
XFILLER_0_18_10 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__1762__A _2200_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_1201_ _2248_/Q _2249_/Q vssd1 vssd1 vccd1 vccd1 _1201_/X sky130_fd_sc_hd__and2_4
X_2181_ _2182_/CLK _2181_/D _1921_/Y vssd1 vssd1 vccd1 vccd1 _2181_/Q sky130_fd_sc_hd__dfrtp_4
X_1132_ _2190_/Q _2098_/Q _1156_/S vssd1 vssd1 vccd1 vccd1 _1132_/X sky130_fd_sc_hd__mux2_1
X_1063_ hold578/X _1097_/A2 _1097_/B1 _1062_/X vssd1 vssd1 vccd1 vccd1 _2313_/D sky130_fd_sc_hd__a22o_1
XFILLER_0_50_41 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_1965_ _2026_/A vssd1 vssd1 vccd1 vccd1 _1965_/Y sky130_fd_sc_hd__inv_2
XFILLER_0_50_85 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__1937__A _1957_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_43_378 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_1896_ _2069_/A vssd1 vssd1 vccd1 vccd1 _1896_/Y sky130_fd_sc_hd__inv_2
XANTENNA__1672__A _2100_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_52_3 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
Xinput209 hold162/X vssd1 vssd1 vccd1 vccd1 hold163/A sky130_fd_sc_hd__clkbuf_1
XANTENNA__1503__B1 _1503_/B1 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_22_518 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_34_356 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__1058__S _1094_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xhold8 hold8/A vssd1 vssd1 vccd1 vccd1 hold8/X sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_38_673 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_1750_ _2188_/Q _1761_/B vssd1 vssd1 vccd1 vccd1 _1750_/X sky130_fd_sc_hd__and2_1
XANTENNA__1757__A _2195_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_37_194 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
Xhold408 hold418/X vssd1 vssd1 vccd1 vccd1 hold408/X sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_20_44 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_1681_ _2109_/Q _1725_/B vssd1 vssd1 vccd1 vccd1 _1681_/X sky130_fd_sc_hd__and2_1
XFILLER_0_52_197 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
Xhold419 _1237_/X vssd1 vssd1 vccd1 vccd1 _2232_/D sky130_fd_sc_hd__dlygate4sd3_1
XTAP_713 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_724 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_702 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_2302_ _2315_/CLK _2302_/D _2041_/Y vssd1 vssd1 vccd1 vccd1 _2302_/Q sky130_fd_sc_hd__dfrtp_1
XTAP_768 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_757 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_746 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_735 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_779 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_2233_ _2238_/CLK _2233_/D _1973_/Y vssd1 vssd1 vccd1 vccd1 _2233_/Q sky130_fd_sc_hd__dfrtp_1
X_2164_ _2164_/CLK hold28/X _1904_/Y vssd1 vssd1 vccd1 vccd1 _2164_/Q sky130_fd_sc_hd__dfrtp_4
X_1115_ hold646/X _1183_/A2 _1183_/B1 _1114_/X vssd1 vssd1 vccd1 vccd1 _2287_/D sky130_fd_sc_hd__a22o_1
XFILLER_0_17_6 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_2095_ _2106_/CLK _2095_/D _1838_/Y vssd1 vssd1 vccd1 vccd1 _2095_/Q sky130_fd_sc_hd__dfrtp_4
X_1046_ _2233_/Q _2141_/Q _1094_/S vssd1 vssd1 vccd1 vccd1 _1046_/X sky130_fd_sc_hd__mux2_1
XFILLER_0_29_673 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_44_632 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__1667__A _2095_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_1948_ _1949_/A vssd1 vssd1 vccd1 vccd1 _1948_/Y sky130_fd_sc_hd__inv_2
X_1879_ _2065_/A vssd1 vssd1 vccd1 vccd1 _1879_/Y sky130_fd_sc_hd__inv_2
XFILLER_0_31_304 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_31_315 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xhold920 _1429_/X vssd1 vssd1 vccd1 vccd1 _2168_/D sky130_fd_sc_hd__dlygate4sd3_1
Xhold931 _2206_/Q vssd1 vssd1 vccd1 vccd1 hold931/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold964 _2089_/Q vssd1 vssd1 vccd1 vccd1 hold964/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold953 _2175_/Q vssd1 vssd1 vccd1 vccd1 hold953/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold942 _2085_/Q vssd1 vssd1 vccd1 vccd1 hold942/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold975 _2182_/Q vssd1 vssd1 vccd1 vccd1 hold975/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold986 _2185_/Q vssd1 vssd1 vccd1 vccd1 hold986/X sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_19_172 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_35_643 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_35_665 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA_hold971_A _2162_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_34_197 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__1516__S _1520_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__1479__C1 hold415/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_output407_A _1725_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_57_278 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_26_654 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_31_76 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_1802_ _2240_/Q _1802_/B vssd1 vssd1 vccd1 vccd1 _1802_/X sky130_fd_sc_hd__and2_1
XFILLER_0_13_326 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_1733_ _2171_/Q _1766_/B vssd1 vssd1 vccd1 vccd1 _1733_/X sky130_fd_sc_hd__and2_2
Xhold205 hold894/X vssd1 vssd1 vccd1 vccd1 hold205/X sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_13_337 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
Xhold216 hold878/X vssd1 vssd1 vccd1 vccd1 hold216/X sky130_fd_sc_hd__dlygate4sd3_1
X_1664_ _2092_/Q _1680_/B vssd1 vssd1 vccd1 vccd1 _1664_/X sky130_fd_sc_hd__and2_1
Xhold238 _1577_/X vssd1 vssd1 vccd1 vccd1 hold238/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold249 _1368_/X vssd1 vssd1 vccd1 vccd1 hold249/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold227 _1331_/X vssd1 vssd1 vccd1 vccd1 hold227/X sky130_fd_sc_hd__buf_1
XFILLER_0_40_178 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__1426__S _1435_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_1595_ input73/X _1619_/A2 _1623_/B1 _2089_/Q _1391_/X vssd1 vssd1 vccd1 vccd1 _1595_/X
+ sky130_fd_sc_hd__a221o_1
XFILLER_0_0_253 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__1182__A1 _2073_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_510 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_521 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_532 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_543 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_565 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_554 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_576 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_2216_ _2217_/CLK _2216_/D _1956_/Y vssd1 vssd1 vccd1 vccd1 _2216_/Q sky130_fd_sc_hd__dfrtp_2
XTAP_587 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_598 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_15_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__1485__A2 _1503_/A2 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_2147_ _2239_/CLK _2147_/D _1890_/Y vssd1 vssd1 vccd1 vccd1 _2147_/Q sky130_fd_sc_hd__dfrtp_2
X_2078_ _2106_/CLK _2078_/D _1821_/Y vssd1 vssd1 vccd1 vccd1 _2078_/Q sky130_fd_sc_hd__dfrtp_4
XFILLER_0_48_234 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_1029_ hold583/X _1057_/A2 _1057_/B1 hold791/X vssd1 vssd1 vccd1 vccd1 _2330_/D sky130_fd_sc_hd__a22o_1
XFILLER_0_36_418 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA_fanout605_A _1949_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_16_197 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_32_657 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_32_668 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_4_592 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xhold750 hold769/X vssd1 vssd1 vccd1 vccd1 hold770/A sky130_fd_sc_hd__buf_1
Xhold761 hold781/X vssd1 vssd1 vccd1 vccd1 hold761/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold772 hold772/A vssd1 vssd1 vccd1 vccd1 hold772/X sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_31_189 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__1336__S hold27/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xhold783 _1197_/C vssd1 vssd1 vccd1 vccd1 hold783/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold794 _2251_/Q vssd1 vssd1 vccd1 vccd1 hold794/X sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA__2021__A _2034_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__1860__A _1949_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_39_223 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_54_215 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_54_259 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_35_473 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_50_432 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_50_421 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_50_454 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__1246__S _1252_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_1380_ input6/X _1529_/A2 _1529_/B1 _2185_/Q hold525/X vssd1 vssd1 vccd1 vccd1 _1380_/X
+ sky130_fd_sc_hd__a221o_1
XANTENNA__1164__A1 _2082_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_clkbuf_leaf_10_wb_clk_i_A clkbuf_1_1__f_wb_clk_i/X vssd1 vssd1 vccd1 vccd1
+ sky130_fd_sc_hd__diode_2
XANTENNA__1770__A _2208_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_2001_ _2008_/A vssd1 vssd1 vccd1 vccd1 _2001_/Y sky130_fd_sc_hd__inv_2
XFILLER_0_45_215 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_45_259 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_5_312 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_26_451 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_53_281 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_41_432 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__1945__A _1949_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_1716_ _2144_/Q _1798_/B vssd1 vssd1 vccd1 vccd1 _1716_/X sky130_fd_sc_hd__and2_1
X_1647_ _2075_/Q _1680_/B vssd1 vssd1 vccd1 vccd1 _1647_/X sky130_fd_sc_hd__and2_1
X_1578_ hold238/X hold956/X _1622_/S vssd1 vssd1 vccd1 vccd1 _2097_/D sky130_fd_sc_hd__mux2_1
XTAP_340 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_351 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xfanout526 hold40/X vssd1 vssd1 vccd1 vccd1 hold26/A sky130_fd_sc_hd__buf_6
Xfanout537 hold79/X vssd1 vssd1 vccd1 vccd1 hold80/A sky130_fd_sc_hd__clkbuf_2
Xfanout548 _1792_/B vssd1 vssd1 vccd1 vccd1 _1761_/B sky130_fd_sc_hd__clkbuf_4
Xfanout559 _1003_/Y vssd1 vssd1 vccd1 vccd1 _1637_/B sky130_fd_sc_hd__buf_4
XTAP_362 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_384 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_373 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__1680__A _2108_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_395 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_fanout555_A _1023_/Y vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XPHY_13 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_24 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_35 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_46 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_57 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_68 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_79 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__2016__A _2034_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__1091__B1 _1097_/B1 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_51_218 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_32_421 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
Xhold580 hold686/X vssd1 vssd1 vccd1 vccd1 hold580/X sky130_fd_sc_hd__clkbuf_2
XANTENNA__1146__A1 _2091_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xhold591 hold724/X vssd1 vssd1 vccd1 vccd1 hold591/X sky130_fd_sc_hd__clkbuf_2
XANTENNA__1749__B _1761_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__1082__A0 _2215_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__1621__A2 _1623_/A2 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_27_248 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_23_421 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__1765__A _2203_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_23_443 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_23_454 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_2_359 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_23_487 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_1501_ _1501_/A1 _1503_/A2 _1503_/B1 _2136_/Q hold325/X vssd1 vssd1 vccd1 vccd1 _1501_/X
+ sky130_fd_sc_hd__a221o_1
X_1432_ hold69/X hold967/X _1435_/S vssd1 vssd1 vccd1 vccd1 _2167_/D sky130_fd_sc_hd__mux2_1
X_1363_ _1362_/X hold947/X _1372_/S vssd1 vssd1 vccd1 vccd1 _2190_/D sky130_fd_sc_hd__mux2_1
X_1294_ hold267/X _2213_/Q _1318_/S vssd1 vssd1 vccd1 vccd1 _1294_/X sky130_fd_sc_hd__mux2_1
XANTENNA__1073__B1 _1095_/B1 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_34_708 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__1675__A _2103_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_14_421 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_14_454 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__1128__A1 _2100_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_192 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_181 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_170 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__1300__A1 _2211_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_49_340 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XANTENNA_hold515_A _1220_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__1064__A0 _2224_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__1603__A2 _1623_/A2 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_45_590 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_58_19 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_20_402 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__1524__S hold80/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_23_11 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_1981_ _1982_/A vssd1 vssd1 vccd1 vccd1 _1981_/Y sky130_fd_sc_hd__inv_2
XFILLER_0_28_557 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_43_505 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_15_218 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_23_295 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_48_63 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_1415_ _1415_/A hold53/X vssd1 vssd1 vccd1 vccd1 hold54/A sky130_fd_sc_hd__and2_1
X_1346_ _1415_/A _1346_/B vssd1 vssd1 vccd1 vccd1 _1346_/X sky130_fd_sc_hd__and2_1
XANTENNA__1530__A1 _2121_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_1277_ _1277_/A _1277_/B vssd1 vssd1 vccd1 vccd1 _1277_/X sky130_fd_sc_hd__and2_1
XFILLER_0_46_332 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_19_535 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_46_365 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XANTENNA__1597__B2 _2088_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_42_571 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
Xoutput471 hold610/X vssd1 vssd1 vccd1 vccd1 la_data_out[56] sky130_fd_sc_hd__buf_12
Xoutput460 hold640/X vssd1 vssd1 vccd1 vccd1 la_data_out[45] sky130_fd_sc_hd__buf_12
XANTENNA_hold298_A _1214_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xoutput482 hold648/X vssd1 vssd1 vccd1 vccd1 la_data_out[67] sky130_fd_sc_hd__buf_12
Xoutput493 hold572/X vssd1 vssd1 vccd1 vccd1 la_data_out[78] sky130_fd_sc_hd__buf_12
XANTENNA__1521__B2 _2126_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__1037__B1 _1095_/B1 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_37_354 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_25_538 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_33_593 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_20_243 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_20_298 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_2180_ _2194_/CLK _2180_/D _1920_/Y vssd1 vssd1 vccd1 vccd1 _2180_/Q sky130_fd_sc_hd__dfrtp_4
X_1200_ hold3/X _2244_/Q _1200_/S vssd1 vssd1 vccd1 vccd1 hold4/A sky130_fd_sc_hd__mux2_1
XANTENNA__1512__A1 _2130_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_1131_ hold598/X _1139_/A2 _1139_/B1 _1130_/X vssd1 vssd1 vccd1 vccd1 _2279_/D sky130_fd_sc_hd__a22o_1
X_1062_ _2225_/Q _2133_/Q _1086_/S vssd1 vssd1 vccd1 vccd1 _1062_/X sky130_fd_sc_hd__mux2_1
XFILLER_0_47_118 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_47_107 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_1964_ _2026_/A vssd1 vssd1 vccd1 vccd1 _1964_/Y sky130_fd_sc_hd__inv_2
XFILLER_0_28_365 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_55_162 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__1579__B2 _2097_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_28_398 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XANTENNA__1429__S _1435_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_43_357 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_43_346 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_1895_ _2069_/A vssd1 vssd1 vccd1 vccd1 _1895_/Y sky130_fd_sc_hd__inv_2
XFILLER_0_3_421 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_11_298 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_45_3 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XANTENNA__1164__S _1188_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__1503__A1 _1503_/A1 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_1329_ input25/X _1197_/D _1541_/B1 _2202_/Q hold254/X vssd1 vssd1 vccd1 vccd1 _1329_/X
+ sky130_fd_sc_hd__a221o_1
XFILLER_0_46_195 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__1863__A _1941_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_30_563 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
Xoutput290 _1766_/X vssd1 vssd1 vccd1 vccd1 data_out[124] sky130_fd_sc_hd__buf_12
Xhold9 hold9/A vssd1 vssd1 vccd1 vccd1 hold9/X sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_57_449 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_37_162 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__1757__B _1792_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_52_121 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_20_23 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__1249__S _1252_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_52_165 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
Xhold409 hold409/A vssd1 vssd1 vccd1 vccd1 _1235_/B sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_20_56 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_1680_ _2108_/Q _1680_/B vssd1 vssd1 vccd1 vccd1 _1680_/X sky130_fd_sc_hd__and2_1
XFILLER_0_0_402 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__1773__A _2211_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_0_424 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_714 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_725 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_703 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_2301_ _2312_/CLK _2301_/D _2040_/Y vssd1 vssd1 vccd1 vccd1 _2301_/Q sky130_fd_sc_hd__dfrtp_1
XTAP_758 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_747 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_736 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_29_65 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_769 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_2232_ _2239_/CLK _2232_/D _1972_/Y vssd1 vssd1 vccd1 vccd1 _2232_/Q sky130_fd_sc_hd__dfrtp_1
X_2163_ _2164_/CLK hold41/X _1903_/Y vssd1 vssd1 vccd1 vccd1 _2163_/Q sky130_fd_sc_hd__dfrtp_4
XFILLER_0_45_53 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_1114_ _2199_/Q _2107_/Q _1178_/S vssd1 vssd1 vccd1 vccd1 _1114_/X sky130_fd_sc_hd__mux2_1
X_2094_ _2106_/CLK _2094_/D _1837_/Y vssd1 vssd1 vccd1 vccd1 _2094_/Q sky130_fd_sc_hd__dfrtp_4
XFILLER_0_48_405 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_1045_ hold650/X _1095_/A2 _1095_/B1 _1044_/X vssd1 vssd1 vccd1 vccd1 _2322_/D sky130_fd_sc_hd__a22o_1
XFILLER_0_48_449 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__1948__A _1949_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_1947_ _1949_/A vssd1 vssd1 vccd1 vccd1 _1947_/Y sky130_fd_sc_hd__inv_2
XFILLER_0_43_165 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_31_327 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_1878_ _2039_/A vssd1 vssd1 vccd1 vccd1 _1878_/Y sky130_fd_sc_hd__inv_2
Xhold921 _2102_/Q vssd1 vssd1 vccd1 vccd1 hold921/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold910 _2143_/Q vssd1 vssd1 vccd1 vccd1 hold910/X sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_12_530 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__1683__A _2111_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xhold932 _2082_/Q vssd1 vssd1 vccd1 vccd1 hold932/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold954 _1408_/X vssd1 vssd1 vccd1 vccd1 _2175_/D sky130_fd_sc_hd__dlygate4sd3_1
Xhold943 _1602_/X vssd1 vssd1 vccd1 vccd1 _2085_/D sky130_fd_sc_hd__dlygate4sd3_1
Xhold987 _2105_/Q vssd1 vssd1 vccd1 vccd1 hold987/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold976 _2203_/Q vssd1 vssd1 vccd1 vccd1 hold976/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold965 _2073_/Q vssd1 vssd1 vccd1 vccd1 hold965/X sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA_fanout585_A _1112_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_39_449 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__1858__A _1949_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_35_622 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA_hold797_A _2113_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_34_154 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_34_187 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA_hold964_A _2089_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_30_382 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_30_393 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__1479__B1 _1503_/B1 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__1532__S hold80/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_15_23 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_57_213 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_15_67 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_45_408 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XANTENNA__1768__A _2206_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_1801_ _2239_/Q _1802_/B vssd1 vssd1 vccd1 vccd1 _1801_/X sky130_fd_sc_hd__and2_1
XFILLER_0_31_11 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_38_460 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_25_110 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_1732_ _2170_/Q _1756_/B vssd1 vssd1 vccd1 vccd1 _1732_/X sky130_fd_sc_hd__and2_1
XFILLER_0_41_625 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_41_603 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_31_88 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_1663_ _2091_/Q _1680_/B vssd1 vssd1 vccd1 vccd1 _1663_/X sky130_fd_sc_hd__and2_1
Xhold206 hold211/X vssd1 vssd1 vccd1 vccd1 hold206/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold217 hold234/X vssd1 vssd1 vccd1 vccd1 hold217/X sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_40_124 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xhold239 hold842/X vssd1 vssd1 vccd1 vccd1 hold239/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold228 _1332_/X vssd1 vssd1 vccd1 vccd1 hold228/X sky130_fd_sc_hd__dlygate4sd3_1
X_1594_ _1593_/X hold964/X _1622_/S vssd1 vssd1 vccd1 vccd1 _2089_/D sky130_fd_sc_hd__mux2_1
XTAP_500 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_511 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_522 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_533 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_0_298 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_544 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_566 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_555 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_2215_ _2217_/CLK _2215_/D _1955_/Y vssd1 vssd1 vccd1 vccd1 _2215_/Q sky130_fd_sc_hd__dfrtp_4
XTAP_577 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_588 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_599 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_56_85 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_2146_ _2224_/CLK _2146_/D _1889_/Y vssd1 vssd1 vccd1 vccd1 _2146_/Q sky130_fd_sc_hd__dfrtp_1
X_2077_ _2182_/CLK _2077_/D _1820_/Y vssd1 vssd1 vccd1 vccd1 _2077_/Q sky130_fd_sc_hd__dfrtp_4
X_1028_ _2242_/Q hold790/X _1094_/S vssd1 vssd1 vccd1 vccd1 _1028_/X sky130_fd_sc_hd__mux2_1
XANTENNA__1678__A _2106_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_29_482 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_8_387 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_8_365 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_44_452 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_32_614 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_12_371 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xhold773 la_data_in[16] vssd1 vssd1 vccd1 vccd1 hold773/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold751 hold751/A vssd1 vssd1 vccd1 vccd1 la_data_out[125] sky130_fd_sc_hd__buf_12
Xhold762 _2154_/Q vssd1 vssd1 vccd1 vccd1 hold762/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold740 hold839/X vssd1 vssd1 vccd1 vccd1 hold740/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold784 _0994_/X vssd1 vssd1 vccd1 vccd1 hold38/A sky130_fd_sc_hd__dlygate4sd3_1
Xhold795 _2302_/Q vssd1 vssd1 vccd1 vccd1 hold795/X sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA__1173__A2 _1183_/A2 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xclkbuf_leaf_18_wb_clk_i clkbuf_1_1__f_wb_clk_i/X vssd1 vssd1 vccd1 vccd1 _2322_/CLK
+ sky130_fd_sc_hd__clkbuf_16
XFILLER_0_35_430 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_50_400 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_23_614 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_35_452 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_35_485 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_22_168 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_22_179 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_30_190 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_2000_ _2008_/A vssd1 vssd1 vccd1 vccd1 _2000_/Y sky130_fd_sc_hd__inv_2
XFILLER_0_26_33 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA_clkbuf_leaf_6_wb_clk_i_A clkbuf_leaf_9_wb_clk_i/A vssd1 vssd1 vccd1 vccd1
+ sky130_fd_sc_hd__diode_2
XFILLER_0_42_43 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_42_32 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_42_65 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_53_293 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_1715_ _2143_/Q _1715_/B vssd1 vssd1 vccd1 vccd1 _1715_/X sky130_fd_sc_hd__and2_1
XFILLER_0_41_466 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_14_669 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_1646_ _2074_/Q _1725_/B vssd1 vssd1 vccd1 vccd1 _1646_/X sky130_fd_sc_hd__and2_1
X_1577_ input83/X _1619_/A2 _1619_/B1 _2098_/Q hold237/X vssd1 vssd1 vccd1 vccd1 _1577_/X
+ sky130_fd_sc_hd__a221o_1
XANTENNA__1961__A _2002_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__1155__A2 _1189_/A2 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xfanout527 _1157_/A2 vssd1 vssd1 vccd1 vccd1 _1189_/A2 sky130_fd_sc_hd__buf_4
XTAP_330 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_341 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xfanout538 _1520_/S vssd1 vssd1 vccd1 vccd1 _1504_/S sky130_fd_sc_hd__buf_6
Xfanout549 _1802_/B vssd1 vssd1 vccd1 vccd1 _1798_/B sky130_fd_sc_hd__clkbuf_4
XTAP_352 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_363 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_385 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_374 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_396 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__1172__S _1188_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_2129_ _2225_/CLK _2129_/D _1872_/Y vssd1 vssd1 vccd1 vccd1 _2129_/Q sky130_fd_sc_hd__dfrtp_2
XPHY_14 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_25 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_36 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_47 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA_fanout548_A _1792_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XPHY_58 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_69 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_49_588 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_32_400 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_32_411 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_32_433 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
Xhold581 hold721/X vssd1 vssd1 vccd1 vccd1 hold581/X sky130_fd_sc_hd__buf_1
XFILLER_0_13_691 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
Xhold570 hold717/X vssd1 vssd1 vccd1 vccd1 hold570/X sky130_fd_sc_hd__clkbuf_2
XANTENNA__1871__A _2002_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xhold592 hold676/X vssd1 vssd1 vccd1 vccd1 hold592/X sky130_fd_sc_hd__dlymetal6s2s_1
XANTENNA_hold927_A _2094_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_27_205 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_55_547 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__1082__A1 _2123_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_12_35 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_35_293 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_11_628 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_23_477 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_23_499 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_1500_ _1499_/X _2136_/Q _1504_/S vssd1 vssd1 vccd1 vccd1 _1500_/X sky130_fd_sc_hd__mux2_1
X_1431_ _1431_/A1 _1569_/A2 _1569_/B1 _2168_/Q hold68/X vssd1 vssd1 vccd1 vccd1 hold69/A
+ sky130_fd_sc_hd__a221o_1
XFILLER_0_10_138 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__2161__GATE_N _1193_/Y vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__1781__A _2219_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_1362_ input13/X _1529_/A2 _1533_/B1 _2191_/Q hold223/X vssd1 vssd1 vccd1 vccd1 _1362_/X
+ sky130_fd_sc_hd__a221o_1
X_1293_ input38/X _1529_/A2 _1529_/B1 _2214_/Q hold266/X vssd1 vssd1 vccd1 vccd1 _1293_/X
+ sky130_fd_sc_hd__a221o_1
Xinput190 hold104/X vssd1 vssd1 vccd1 vccd1 hold105/A sky130_fd_sc_hd__clkbuf_1
XFILLER_0_46_514 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__1021__A hold38/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_18_205 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_46_536 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__1956__A _1957_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_14_477 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_1629_ input75/X _1637_/B _1635_/C _2072_/Q hold31/X vssd1 vssd1 vccd1 vccd1 hold32/A
+ sky130_fd_sc_hd__a221o_1
XANTENNA__1691__A _2119_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_160 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_193 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_182 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_171 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_49_352 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__2027__A _2034_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_37_503 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_37_536 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_45_580 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_32_230 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_20_414 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__1119__A2 _1189_/A2 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__1540__S hold80/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_1980_ _1982_/A vssd1 vssd1 vccd1 vccd1 _1980_/Y sky130_fd_sc_hd__inv_2
XFILLER_0_28_525 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_55_311 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_28_536 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__1776__A _2214_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_43_517 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_11_447 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_48_75 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_1414_ _1413_/X _2173_/Q hold27/X vssd1 vssd1 vccd1 vccd1 _1414_/X sky130_fd_sc_hd__mux2_1
X_1345_ _1344_/X hold935/X _1435_/S vssd1 vssd1 vccd1 vccd1 _1345_/X sky130_fd_sc_hd__mux2_1
XFILLER_0_3_66 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_1276_ hold341/X hold974/X _1318_/S vssd1 vssd1 vccd1 vccd1 _2219_/D sky130_fd_sc_hd__mux2_1
XANTENNA__1294__A1 _2213_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_19_503 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_46_377 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_46_344 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XANTENNA__1686__A _2114_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_14_241 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_42_594 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xoutput461 hold608/X vssd1 vssd1 vccd1 vccd1 la_data_out[46] sky130_fd_sc_hd__buf_12
Xoutput450 hold625/X vssd1 vssd1 vccd1 vccd1 la_data_out[35] sky130_fd_sc_hd__buf_12
Xoutput483 hold649/X vssd1 vssd1 vccd1 vccd1 la_data_out[68] sky130_fd_sc_hd__buf_12
Xoutput472 hold597/X vssd1 vssd1 vccd1 vccd1 la_data_out[57] sky130_fd_sc_hd__buf_12
Xoutput494 hold586/X vssd1 vssd1 vccd1 vccd1 la_data_out[79] sky130_fd_sc_hd__buf_12
XANTENNA__1521__A2 _1527_/A2 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__1285__A1 _2216_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_37_311 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_37_366 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_25_528 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_37_399 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_1130_ _2191_/Q _2099_/Q _1156_/S vssd1 vssd1 vccd1 vccd1 _1130_/X sky130_fd_sc_hd__mux2_1
XANTENNA__1270__S _1318_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_1061_ hold644/X _1095_/A2 _1095_/B1 _1060_/X vssd1 vssd1 vccd1 vccd1 _2314_/D sky130_fd_sc_hd__a22o_1
XFILLER_0_34_66 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_56_642 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_1963_ _2002_/A vssd1 vssd1 vccd1 vccd1 _1963_/Y sky130_fd_sc_hd__inv_2
XFILLER_0_28_344 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_28_355 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_50_65 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_43_325 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_1894_ _1949_/A vssd1 vssd1 vccd1 vccd1 _1894_/Y sky130_fd_sc_hd__inv_2
XFILLER_0_51_391 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__1503__A2 _1503_/A2 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_38_3 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_1328_ _1349_/A _1328_/B vssd1 vssd1 vccd1 vccd1 _1328_/X sky130_fd_sc_hd__and2_1
X_1259_ _1277_/A _1259_/B vssd1 vssd1 vccd1 vccd1 _1259_/X sky130_fd_sc_hd__and2_1
XANTENNA__1180__S _1188_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__1267__A1 _2222_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_38_108 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_46_141 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_30_531 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_30_553 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
Xoutput280 _1757_/X vssd1 vssd1 vccd1 vccd1 data_out[115] sky130_fd_sc_hd__buf_12
XANTENNA__2040__A _2065_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xoutput291 _1767_/X vssd1 vssd1 vccd1 vccd1 data_out[125] sky130_fd_sc_hd__buf_12
XANTENNA__1090__S _1094_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_38_653 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_38_664 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_38_686 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_40_306 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_40_317 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_715 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_704 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_29_44 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_2300_ _2300_/CLK _2300_/D _2039_/Y vssd1 vssd1 vccd1 vccd1 _2300_/Q sky130_fd_sc_hd__dfrtp_1
XTAP_759 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_748 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_737 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_726 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_2231_ _2239_/CLK _2231_/D _1971_/Y vssd1 vssd1 vccd1 vccd1 _2231_/Q sky130_fd_sc_hd__dfrtp_1
X_2162_ _2173_/CLK _2162_/D _1902_/Y vssd1 vssd1 vccd1 vccd1 _2162_/Q sky130_fd_sc_hd__dfrtp_4
XANTENNA__1497__A1 _1497_/A1 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_1113_ hold584/X _1183_/A2 _1183_/B1 _1112_/X vssd1 vssd1 vccd1 vccd1 _2288_/D sky130_fd_sc_hd__a22o_1
X_2093_ _2106_/CLK _2093_/D _1836_/Y vssd1 vssd1 vccd1 vccd1 _2093_/Q sky130_fd_sc_hd__dfrtp_4
X_1044_ _2234_/Q _2142_/Q _1086_/S vssd1 vssd1 vccd1 vccd1 _1044_/X sky130_fd_sc_hd__mux2_1
XFILLER_0_28_152 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_44_645 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_43_111 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_1946_ _1949_/A vssd1 vssd1 vccd1 vccd1 _1946_/Y sky130_fd_sc_hd__inv_2
XANTENNA__1964__A _2026_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_1877_ _2039_/A vssd1 vssd1 vccd1 vccd1 _1877_/Y sky130_fd_sc_hd__inv_2
Xhold922 _2179_/Q vssd1 vssd1 vccd1 vccd1 hold922/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold900 la_data_in[10] vssd1 vssd1 vccd1 vccd1 hold900/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold911 _2276_/Q vssd1 vssd1 vccd1 vccd1 hold911/X sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_24_380 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_24_391 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xhold944 _2192_/Q vssd1 vssd1 vccd1 vccd1 hold944/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold955 _2183_/Q vssd1 vssd1 vccd1 vccd1 hold955/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold933 _2103_/Q vssd1 vssd1 vccd1 vccd1 hold933/X sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA__1683__B _1725_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xhold966 _2181_/Q vssd1 vssd1 vccd1 vccd1 hold966/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold977 _2169_/Q vssd1 vssd1 vccd1 vccd1 hold977/X sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA__1185__B1 _1189_/B1 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xhold988 _2172_/Q vssd1 vssd1 vccd1 vccd1 hold988/X sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA_fanout578_A _1529_/B1 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__1204__A hold38/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_47_472 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_19_152 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__2035__A _2065_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__1874__A _2002_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_35_689 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__1176__A0 _2168_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_15_391 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA_hold957_A _2218_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__1479__A1 _1479_/A1 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__1479__B2 _2147_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_15_57 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_57_225 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__1100__A0 _2206_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_1800_ _2238_/Q _1802_/B vssd1 vssd1 vccd1 vccd1 _1800_/X sky130_fd_sc_hd__and2_1
XFILLER_0_26_645 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_31_45 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_1731_ _2169_/Q _1756_/B vssd1 vssd1 vccd1 vccd1 _1731_/X sky130_fd_sc_hd__and2_1
XANTENNA__1784__A _2222_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_1662_ _2090_/Q _1680_/B vssd1 vssd1 vccd1 vccd1 _1662_/X sky130_fd_sc_hd__and2_1
Xhold207 hold207/A vssd1 vssd1 vccd1 vccd1 _1370_/B sky130_fd_sc_hd__dlygate4sd3_1
Xhold218 hold218/A vssd1 vssd1 vccd1 vccd1 _1406_/B sky130_fd_sc_hd__dlygate4sd3_1
Xhold229 hold240/X vssd1 vssd1 vccd1 vccd1 hold229/X sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_40_136 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_1593_ input74/X _1619_/A2 _1623_/B1 _2090_/Q _1388_/X vssd1 vssd1 vccd1 vccd1 _1593_/X
+ sky130_fd_sc_hd__a221o_1
XANTENNA__1167__B1 _1183_/B1 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_501 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_512 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_523 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_534 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__1008__B _1811_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_545 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_567 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_556 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_2214_ _2219_/CLK _2214_/D _1954_/Y vssd1 vssd1 vccd1 vccd1 _2214_/Q sky130_fd_sc_hd__dfrtp_4
XTAP_578 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_589 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_2145_ _2224_/CLK _2145_/D _1888_/Y vssd1 vssd1 vccd1 vccd1 _2145_/Q sky130_fd_sc_hd__dfrtp_2
X_2076_ _2168_/CLK hold82/X _1819_/Y vssd1 vssd1 vccd1 vccd1 _2076_/Q sky130_fd_sc_hd__dfrtp_4
XFILLER_0_48_214 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_1027_ hold88/X _1198_/B _1198_/C vssd1 vssd1 vccd1 vccd1 _1027_/Y sky130_fd_sc_hd__nand3_1
XANTENNA__1959__A _2002_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_1929_ _1941_/A vssd1 vssd1 vccd1 vccd1 _1929_/Y sky130_fd_sc_hd__inv_2
XFILLER_0_44_464 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_32_604 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_44_497 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_31_125 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_32_637 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
Xhold730 hold897/X vssd1 vssd1 vccd1 vccd1 hold730/X sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_31_169 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
Xhold752 hold771/X vssd1 vssd1 vccd1 vccd1 hold772/A sky130_fd_sc_hd__buf_1
Xhold741 hold911/X vssd1 vssd1 vccd1 vccd1 hold741/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold763 _2291_/Q vssd1 vssd1 vccd1 vccd1 hold763/X sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA__1158__A0 _2177_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xhold774 _1600_/X vssd1 vssd1 vccd1 vccd1 _2086_/D sky130_fd_sc_hd__dlygate4sd3_1
Xhold785 la_data_in[92] vssd1 vssd1 vccd1 vccd1 hold785/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold796 _2288_/Q vssd1 vssd1 vccd1 vccd1 hold796/X sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA__1869__A _2002_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_39_225 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_27_409 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_39_247 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_54_239 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_35_442 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_23_637 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_35_497 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_10_309 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__1149__B1 _1183_/B1 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xhold90 hold90/A vssd1 vssd1 vccd1 vccd1 hold90/X sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA__1779__A _2217_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_26_475 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_1714_ _2142_/Q _1756_/B vssd1 vssd1 vccd1 vccd1 _1714_/X sky130_fd_sc_hd__and2_1
XFILLER_0_6_33 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_6_11 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_1645_ _2073_/Q _1725_/B vssd1 vssd1 vccd1 vccd1 _1645_/X sky130_fd_sc_hd__and2_1
X_1576_ hold224/X hold962/X _1622_/S vssd1 vssd1 vccd1 vccd1 _2098_/D sky130_fd_sc_hd__mux2_1
Xfanout539 hold79/X vssd1 vssd1 vccd1 vccd1 _1520_/S sky130_fd_sc_hd__clkbuf_8
Xfanout528 _1157_/A2 vssd1 vssd1 vccd1 vccd1 _1139_/A2 sky130_fd_sc_hd__buf_2
XFILLER_0_6_99 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_320 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_331 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_342 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_353 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_364 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_375 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_386 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_397 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_20_3 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_49_501 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_2128_ _2256_/CLK _2128_/D _1871_/Y vssd1 vssd1 vccd1 vccd1 _2128_/Q sky130_fd_sc_hd__dfrtp_2
XPHY_15 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_2059_ _2069_/A vssd1 vssd1 vccd1 vccd1 _2059_/Y sky130_fd_sc_hd__inv_2
XPHY_26 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_37 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__1689__A _2117_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_49_556 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_9_620 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XPHY_48 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_59 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_8_130 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__1615__B2 _2079_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__1091__A2 _1097_/A2 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout610_A _2026_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_17_442 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_44_294 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_20_607 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_20_629 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xhold560 _0965_/X vssd1 vssd1 vccd1 vccd1 _0966_/D sky130_fd_sc_hd__dlygate4sd3_1
Xhold571 hold707/X vssd1 vssd1 vccd1 vccd1 hold571/X sky130_fd_sc_hd__dlymetal6s2s_1
Xhold582 _1466_/X vssd1 vssd1 vccd1 vccd1 _2152_/D sky130_fd_sc_hd__dlygate4sd3_1
Xhold593 hold667/X vssd1 vssd1 vccd1 vccd1 hold593/X sky130_fd_sc_hd__dlymetal6s2s_1
XFILLER_0_59_309 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_12_58 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__1538__S hold80/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_2_306 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_2_328 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_50_253 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_10_128 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_1430_ _1445_/A hold67/X vssd1 vssd1 vccd1 vccd1 hold68/A sky130_fd_sc_hd__and2_1
X_1361_ _1415_/A _1361_/B vssd1 vssd1 vccd1 vccd1 _1361_/X sky130_fd_sc_hd__and2_1
XANTENNA__1273__S _1318_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_37_33 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_1292_ _1310_/A _1292_/B vssd1 vssd1 vccd1 vccd1 _1292_/X sky130_fd_sc_hd__and2_1
XFILLER_0_37_55 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xinput180 hold125/X vssd1 vssd1 vccd1 vccd1 hold126/A sky130_fd_sc_hd__clkbuf_1
Xinput191 hold134/X vssd1 vssd1 vccd1 vccd1 hold135/A sky130_fd_sc_hd__buf_1
XFILLER_0_53_76 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
Xclkbuf_leaf_3_wb_clk_i clkbuf_leaf_9_wb_clk_i/A vssd1 vssd1 vccd1 vccd1 _2106_/CLK
+ sky130_fd_sc_hd__clkbuf_16
XANTENNA__1073__A2 _1095_/A2 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_26_272 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_14_445 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_26_294 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__1230__C1 hold348/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_41_275 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_41_253 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XANTENNA__1972__A _1979_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_1628_ hold18/X _2072_/Q _1632_/S vssd1 vssd1 vccd1 vccd1 hold19/A sky130_fd_sc_hd__mux2_1
XFILLER_0_10_651 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__1691__B _1724_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_1559_ input93/X _1623_/A2 _1623_/B1 _2107_/Q hold344/X vssd1 vssd1 vccd1 vccd1 _1559_/X
+ sky130_fd_sc_hd__a221o_1
XTAP_150 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_183 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_172 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_161 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_194 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_fanout560_A _1003_/Y vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_37_559 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_24_209 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_33_710 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__2043__A _2065_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_32_242 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__1221__C1 hold515/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_32_253 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__1882__A _1979_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xhold390 hold390/A vssd1 vssd1 vccd1 vccd1 _1280_/B sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA__1055__A2 _1095_/A2 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_43_529 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__1515__B1 _1519_/B1 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_1413_ _1413_/A1 _1198_/A _1545_/B1 _2174_/Q hold156/X vssd1 vssd1 vccd1 vccd1 _1413_/X
+ sky130_fd_sc_hd__a221o_1
X_1344_ input19/X _1533_/A2 _1533_/B1 _2197_/Q hold136/X vssd1 vssd1 vccd1 vccd1 _1344_/X
+ sky130_fd_sc_hd__a221o_1
X_1275_ input44/X _1529_/A2 _1529_/B1 _2220_/Q hold340/X vssd1 vssd1 vccd1 vccd1 _1275_/X
+ sky130_fd_sc_hd__a221o_1
XFILLER_0_59_673 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__1967__A _1979_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_46_356 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__1686__B _1725_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_27_581 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_6_475 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_42_562 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_14_253 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_30_713 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_42_584 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xoutput440 hold702/X vssd1 vssd1 vccd1 vccd1 hold703/A sky130_fd_sc_hd__buf_6
Xoutput451 hold628/X vssd1 vssd1 vccd1 vccd1 la_data_out[36] sky130_fd_sc_hd__buf_12
Xoutput462 hold606/X vssd1 vssd1 vccd1 vccd1 la_data_out[47] sky130_fd_sc_hd__buf_12
Xoutput495 hold579/X vssd1 vssd1 vccd1 vccd1 la_data_out[80] sky130_fd_sc_hd__buf_12
Xoutput473 hold600/X vssd1 vssd1 vccd1 vccd1 la_data_out[58] sky130_fd_sc_hd__buf_12
Xoutput484 hold646/X vssd1 vssd1 vccd1 vccd1 la_data_out[69] sky130_fd_sc_hd__buf_12
XANTENNA__1037__A2 _1095_/A2 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_37_301 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__1877__A _2039_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__1088__S _1112_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_52_337 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XANTENNA_hold987_A _2105_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_21_702 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_20_256 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_18_13 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_1060_ _2226_/Q _2134_/Q _1086_/S vssd1 vssd1 vccd1 vccd1 _1060_/X sky130_fd_sc_hd__mux2_1
XFILLER_0_34_23 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_34_45 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_28_312 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_1962_ _2002_/A vssd1 vssd1 vccd1 vccd1 _1962_/Y sky130_fd_sc_hd__inv_2
XFILLER_0_56_698 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_43_304 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_1893_ _1982_/A vssd1 vssd1 vccd1 vccd1 _1893_/Y sky130_fd_sc_hd__inv_2
XFILLER_0_50_77 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_43_337 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_12_713 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_51_381 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_1327_ _1326_/X _2202_/Q hold27/X vssd1 vssd1 vccd1 vccd1 _1327_/X sky130_fd_sc_hd__mux2_1
X_1258_ _1257_/X _2225_/Q hold26/X vssd1 vssd1 vccd1 vccd1 _1258_/X sky130_fd_sc_hd__mux2_1
X_1189_ hold605/X _1189_/A2 _1189_/B1 _1188_/X vssd1 vssd1 vccd1 vccd1 _2250_/D sky130_fd_sc_hd__a22o_1
XANTENNA__1697__A _2125_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_19_301 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA_fanout523_A hold26/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_46_164 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_19_378 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xoutput270 _1748_/X vssd1 vssd1 vccd1 vccd1 data_out[106] sky130_fd_sc_hd__buf_12
XFILLER_0_30_587 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xoutput292 _1768_/X vssd1 vssd1 vccd1 vccd1 data_out[126] sky130_fd_sc_hd__buf_12
Xoutput281 _1758_/X vssd1 vssd1 vccd1 vccd1 data_out[116] sky130_fd_sc_hd__buf_12
XANTENNA__1400__A _1415_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_25_337 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_52_178 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_20_47 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_33_370 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_40_329 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_716 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_705 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_749 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_738 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_727 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_29_78 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_2230_ _2239_/CLK _2230_/D _1970_/Y vssd1 vssd1 vccd1 vccd1 _2230_/Q sky130_fd_sc_hd__dfrtp_1
XFILLER_0_45_22 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_2161_ _2161_/D _1193_/Y vssd1 vssd1 vccd1 vccd1 _2161_/Q sky130_fd_sc_hd__dlxtn_1
X_2092_ _2182_/CLK _2092_/D _1835_/Y vssd1 vssd1 vccd1 vccd1 _2092_/Q sky130_fd_sc_hd__dfrtp_4
X_1112_ _2200_/Q _2108_/Q _1112_/S vssd1 vssd1 vccd1 vccd1 _1112_/X sky130_fd_sc_hd__mux2_1
X_1043_ hold596/X _1057_/A2 _1057_/B1 _1042_/X vssd1 vssd1 vccd1 vccd1 _2323_/D sky130_fd_sc_hd__a22o_1
XFILLER_0_17_9 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_48_429 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_29_610 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__1310__A _1310_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_29_643 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_29_654 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_1945_ _1949_/A vssd1 vssd1 vccd1 vccd1 _1945_/Y sky130_fd_sc_hd__inv_2
XFILLER_0_44_635 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_28_197 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_43_156 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_31_318 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_1876_ _2002_/A vssd1 vssd1 vccd1 vccd1 _1876_/Y sky130_fd_sc_hd__inv_2
Xhold912 la_data_in[35] vssd1 vssd1 vccd1 vccd1 hold912/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold901 _1417_/X vssd1 vssd1 vccd1 vccd1 _2172_/D sky130_fd_sc_hd__dlygate4sd3_1
Xhold934 _1566_/X vssd1 vssd1 vccd1 vccd1 _2103_/D sky130_fd_sc_hd__dlygate4sd3_1
Xhold945 _2127_/Q vssd1 vssd1 vccd1 vccd1 hold945/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold923 _2177_/Q vssd1 vssd1 vccd1 vccd1 hold923/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold978 _2195_/Q vssd1 vssd1 vccd1 vccd1 hold978/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold956 _2097_/Q vssd1 vssd1 vccd1 vccd1 hold956/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold967 _2167_/Q vssd1 vssd1 vccd1 vccd1 hold967/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold989 _2111_/Q vssd1 vssd1 vccd1 vccd1 hold989/X sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_50_3 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_19_164 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_22_307 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__2051__A _2065_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__1176__A1 _2076_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__1890__A _1979_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__1479__A2 _1503_/A2 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__1100__A1 _2114_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_26_613 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_31_57 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_1730_ _2168_/Q _1761_/B vssd1 vssd1 vccd1 vccd1 _1730_/X sky130_fd_sc_hd__and2_1
XFILLER_0_25_167 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_31_79 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_1661_ _2089_/Q _1677_/B vssd1 vssd1 vccd1 vccd1 _1661_/X sky130_fd_sc_hd__and2_1
Xhold208 _1370_/X vssd1 vssd1 vccd1 vccd1 hold208/X sky130_fd_sc_hd__dlymetal6s2s_1
XANTENNA__1276__S _1318_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xhold219 _1406_/X vssd1 vssd1 vccd1 vccd1 hold219/X sky130_fd_sc_hd__buf_1
X_1592_ _1591_/X hold980/X _1622_/S vssd1 vssd1 vccd1 vccd1 _2090_/D sky130_fd_sc_hd__mux2_1
XFILLER_0_21_373 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_502 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_513 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_524 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_56_21 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_535 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_557 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_546 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_568 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_579 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_2213_ _2219_/CLK _2213_/D _1953_/Y vssd1 vssd1 vccd1 vccd1 _2213_/Q sky130_fd_sc_hd__dfrtp_4
X_2144_ _2238_/CLK _2144_/D _1887_/Y vssd1 vssd1 vccd1 vccd1 _2144_/Q sky130_fd_sc_hd__dfrtp_1
X_2075_ _2106_/CLK _2075_/D _1818_/Y vssd1 vssd1 vccd1 vccd1 _2075_/Q sky130_fd_sc_hd__dfrtp_4
X_1026_ hold88/X _1198_/B _1198_/C vssd1 vssd1 vccd1 vccd1 _1038_/S sky130_fd_sc_hd__and3_4
XFILLER_0_48_259 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_44_421 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__1975__A _1979_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_1928_ _1941_/A vssd1 vssd1 vccd1 vccd1 _1928_/Y sky130_fd_sc_hd__inv_2
XANTENNA__1694__B _1715_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__1186__S _1188_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_1859_ _1949_/A vssd1 vssd1 vccd1 vccd1 _1859_/Y sky130_fd_sc_hd__inv_2
Xhold720 hold856/X vssd1 vssd1 vccd1 vccd1 hold720/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold742 hold764/X vssd1 vssd1 vccd1 vccd1 hold742/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold753 hold753/A vssd1 vssd1 vccd1 vccd1 la_data_out[124] sky130_fd_sc_hd__buf_12
Xhold731 hold850/X vssd1 vssd1 vccd1 vccd1 hold731/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold764 _2272_/Q vssd1 vssd1 vccd1 vccd1 hold764/X sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA__1158__A1 _2085_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xhold775 _2178_/Q vssd1 vssd1 vccd1 vccd1 hold775/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold797 _2113_/Q vssd1 vssd1 vccd1 vccd1 hold797/X sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA_fanout590_A _1038_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xhold786 _2109_/Q vssd1 vssd1 vccd1 vccd1 hold786/X sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA__2046__A _2065_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__1094__A0 _2209_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__1885__A _2039_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_47_292 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XANTENNA__1096__S _1112_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_50_457 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_22_137 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_31_671 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xhold91 hold91/A vssd1 vssd1 vccd1 vccd1 hold91/X sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA__1321__A1 _2204_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xhold80 hold80/A vssd1 vssd1 vccd1 vccd1 hold80/X sky130_fd_sc_hd__buf_6
XANTENNA_output405_A _1723_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__1085__B1 _1095_/B1 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_26_421 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_38_292 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_53_251 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_5_337 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_53_262 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_1713_ _2141_/Q _1756_/B vssd1 vssd1 vccd1 vccd1 _1713_/X sky130_fd_sc_hd__and2_1
XFILLER_0_41_446 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_1644_ _2072_/Q _1725_/B vssd1 vssd1 vccd1 vccd1 _1644_/X sky130_fd_sc_hd__and2_1
X_1575_ input84/X _1619_/A2 _1619_/B1 _2099_/Q hold223/X vssd1 vssd1 vccd1 vccd1 _1575_/X
+ sky130_fd_sc_hd__a221o_1
XFILLER_0_21_181 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_310 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_321 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_332 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xfanout529 _1157_/A2 vssd1 vssd1 vccd1 vccd1 _1183_/A2 sky130_fd_sc_hd__buf_4
XTAP_343 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_354 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_365 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_376 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_387 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_398 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__1312__A1 _2207_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_2127_ _2219_/CLK _2127_/D _1870_/Y vssd1 vssd1 vccd1 vccd1 _2127_/Q sky130_fd_sc_hd__dfrtp_4
X_2058_ _2069_/A vssd1 vssd1 vccd1 vccd1 _2058_/Y sky130_fd_sc_hd__inv_2
XPHY_16 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_38 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__1689__B _1724_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__1076__A0 _2218_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_1009_ hold561/X _0971_/X _1810_/C vssd1 vssd1 vccd1 vccd1 _1009_/X sky130_fd_sc_hd__a21o_1
XPHY_49 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__1615__A2 _1623_/A2 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_29_281 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA_fanout603_A _1957_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_17_498 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xhold550 hold760/X vssd1 vssd1 vccd1 vccd1 _2245_/D sky130_fd_sc_hd__dlygate4sd3_1
Xhold561 _1455_/B vssd1 vssd1 vccd1 vccd1 hold561/X sky130_fd_sc_hd__buf_1
Xhold572 hold689/X vssd1 vssd1 vccd1 vccd1 hold572/X sky130_fd_sc_hd__clkbuf_2
Xhold594 hold698/X vssd1 vssd1 vccd1 vccd1 hold594/X sky130_fd_sc_hd__buf_1
Xhold583 hold665/X vssd1 vssd1 vccd1 vccd1 hold583/X sky130_fd_sc_hd__buf_1
XANTENNA__1551__B2 _2111_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__1303__A1 _2210_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__1067__B1 _1095_/B1 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_50_243 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_23_457 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_50_276 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_1360_ _1359_/X _2191_/Q _1372_/S vssd1 vssd1 vccd1 vccd1 _1360_/X sky130_fd_sc_hd__mux2_1
XANTENNA__1542__A1 _2115_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_1291_ hold286/X _2214_/Q _1318_/S vssd1 vssd1 vccd1 vccd1 _1291_/X sky130_fd_sc_hd__mux2_1
Xinput181 hold206/X vssd1 vssd1 vccd1 vccd1 hold207/A sky130_fd_sc_hd__buf_1
Xinput170 hold130/X vssd1 vssd1 vccd1 vccd1 hold131/A sky130_fd_sc_hd__clkbuf_1
Xinput192 hold367/X vssd1 vssd1 vccd1 vccd1 hold368/A sky130_fd_sc_hd__clkbuf_1
XFILLER_0_53_88 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XANTENNA__1230__B1 _1503_/B1 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_41_265 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_1627_ input86/X _1637_/B _1635_/C _2073_/Q hold17/X vssd1 vssd1 vccd1 vccd1 hold18/A
+ sky130_fd_sc_hd__a221o_1
XTAP_140 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__1533__B2 _2120_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_1558_ _1557_/X _2107_/Q hold81/X vssd1 vssd1 vccd1 vccd1 _1558_/X sky130_fd_sc_hd__mux2_1
X_1489_ _1489_/A1 _1503_/A2 _1503_/B1 _2142_/Q hold384/X vssd1 vssd1 vccd1 vccd1 _1489_/X
+ sky130_fd_sc_hd__a221o_1
XTAP_184 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_173 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_151 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_162 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_195 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_fanout553_A _1157_/B1 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_49_365 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__1049__B1 _1095_/B1 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_37_505 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_17_251 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_17_262 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_17_284 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__1221__B1 _1503_/B1 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_20_405 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xhold380 _1497_/X vssd1 vssd1 vccd1 vccd1 hold380/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold391 _1280_/X vssd1 vssd1 vccd1 vccd1 hold391/X sky130_fd_sc_hd__buf_1
XANTENNA_hold932_A _2082_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__1403__A _1415_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_28_516 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_55_335 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__1460__B1 _1541_/B1 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_36_571 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_2_104 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_23_298 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__1792__B _1792_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_1412_ _1415_/A _1412_/B vssd1 vssd1 vccd1 vccd1 _1412_/X sky130_fd_sc_hd__and2_1
XANTENNA__1515__A1 _1515_/A1 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_1343_ _1415_/A _1343_/B vssd1 vssd1 vccd1 vccd1 _1343_/X sky130_fd_sc_hd__and2_1
X_1274_ _1277_/A _1274_/B vssd1 vssd1 vccd1 vccd1 _1274_/X sky130_fd_sc_hd__and2_1
XFILLER_0_3_57 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_19_538 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_6_421 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_54_390 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_0989_ _0992_/A _0992_/B vssd1 vssd1 vccd1 vccd1 _1014_/D sky130_fd_sc_hd__and2_1
XFILLER_0_27_593 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_14_265 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
Xoutput441 hold768/X vssd1 vssd1 vccd1 vccd1 hold749/A sky130_fd_sc_hd__buf_6
Xoutput430 hold595/X vssd1 vssd1 vccd1 vccd1 la_data_out[103] sky130_fd_sc_hd__buf_12
Xoutput452 hold604/X vssd1 vssd1 vccd1 vccd1 la_data_out[37] sky130_fd_sc_hd__buf_12
Xoutput485 hold584/X vssd1 vssd1 vccd1 vccd1 la_data_out[70] sky130_fd_sc_hd__buf_12
Xoutput474 hold614/X vssd1 vssd1 vccd1 vccd1 la_data_out[59] sky130_fd_sc_hd__buf_12
Xoutput463 hold567/X vssd1 vssd1 vccd1 vccd1 la_data_out[48] sky130_fd_sc_hd__buf_12
Xoutput496 hold574/X vssd1 vssd1 vccd1 vccd1 la_data_out[81] sky130_fd_sc_hd__buf_12
XFILLER_0_49_151 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_49_140 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xclkbuf_1_1__f_wb_clk_i clkbuf_0_wb_clk_i/X vssd1 vssd1 vccd1 vccd1 clkbuf_1_1__f_wb_clk_i/X
+ sky130_fd_sc_hd__clkbuf_16
XFILLER_0_9_270 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_18_571 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_52_349 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_33_585 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_18_47 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__1279__S _1318_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_1961_ _2002_/A vssd1 vssd1 vccd1 vccd1 _1961_/Y sky130_fd_sc_hd__inv_2
XFILLER_0_55_165 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_1892_ _1982_/A vssd1 vssd1 vccd1 vccd1 _1892_/Y sky130_fd_sc_hd__inv_2
XFILLER_0_51_393 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_1326_ input26/X _1197_/D _1541_/B1 _2203_/Q hold191/X vssd1 vssd1 vccd1 vccd1 _1326_/X
+ sky130_fd_sc_hd__a221o_1
X_1257_ input51/X _1519_/A2 _1519_/B1 _2226_/Q hold475/X vssd1 vssd1 vccd1 vccd1 _1257_/X
+ sky130_fd_sc_hd__a221o_1
X_1188_ hold971/X _2070_/Q _1188_/S vssd1 vssd1 vccd1 vccd1 _1188_/X sky130_fd_sc_hd__mux2_1
XANTENNA__1978__A _2039_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__1697__B _1715_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_46_121 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_46_110 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_19_335 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_19_346 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_46_176 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_6_251 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_27_390 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_42_393 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
Xoutput271 _1749_/X vssd1 vssd1 vccd1 vccd1 data_out[107] sky130_fd_sc_hd__buf_12
XFILLER_0_30_599 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
Xoutput282 _1759_/X vssd1 vssd1 vccd1 vccd1 data_out[117] sky130_fd_sc_hd__buf_12
Xoutput293 _1769_/X vssd1 vssd1 vccd1 vccd1 data_out[127] sky130_fd_sc_hd__buf_12
XFILLER_0_10_290 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__1888__A _2039_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_38_677 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_52_124 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_20_15 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_25_349 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_20_37 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_20_59 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_21_500 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_33_393 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_706 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_739 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_717 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_728 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_29_57 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_2160_ _2251_/CLK _2160_/D _1901_/Y vssd1 vssd1 vccd1 vccd1 _2160_/Q sky130_fd_sc_hd__dfrtp_1
X_2091_ _2182_/CLK _2091_/D _1834_/Y vssd1 vssd1 vccd1 vccd1 _2091_/Q sky130_fd_sc_hd__dfrtp_4
X_1111_ hold585/X _1139_/A2 _1139_/B1 _1110_/X vssd1 vssd1 vccd1 vccd1 _2289_/D sky130_fd_sc_hd__a22o_1
X_1042_ _2235_/Q _2143_/Q _1094_/S vssd1 vssd1 vccd1 vccd1 _1042_/X sky130_fd_sc_hd__mux2_1
XFILLER_0_48_408 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_48_419 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_28_110 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_56_474 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_44_625 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_1944_ _1949_/A vssd1 vssd1 vccd1 vccd1 _1944_/Y sky130_fd_sc_hd__inv_2
X_1875_ _2002_/A vssd1 vssd1 vccd1 vccd1 _1875_/Y sky130_fd_sc_hd__inv_2
Xhold913 _1342_/X vssd1 vssd1 vccd1 vccd1 _2197_/D sky130_fd_sc_hd__dlygate4sd3_1
Xhold902 la_data_in[38] vssd1 vssd1 vccd1 vccd1 hold902/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold924 _2223_/Q vssd1 vssd1 vccd1 vccd1 hold924/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold935 _2196_/Q vssd1 vssd1 vccd1 vccd1 hold935/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold946 _1518_/X vssd1 vssd1 vccd1 vccd1 _2127_/D sky130_fd_sc_hd__dlygate4sd3_1
Xhold957 _2218_/Q vssd1 vssd1 vccd1 vccd1 hold957/X sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA__1185__A2 _1189_/A2 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xhold968 _2199_/Q vssd1 vssd1 vccd1 vccd1 hold968/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold979 _2166_/Q vssd1 vssd1 vccd1 vccd1 hold979/X sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_43_3 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XANTENNA__1472__S _1504_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_2289_ _2291_/CLK _2289_/D _2028_/Y vssd1 vssd1 vccd1 vccd1 _2289_/Q sky130_fd_sc_hd__dfrtp_1
X_1309_ hold60/X _2208_/Q _1318_/S vssd1 vssd1 vccd1 vccd1 hold61/A sky130_fd_sc_hd__mux2_1
XFILLER_0_35_614 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_42_190 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_15_393 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XANTENNA__1581__C1 hold208/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_30_385 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_15_15 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_38_463 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_25_113 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_26_658 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_1660_ _2088_/Q _1677_/B vssd1 vssd1 vccd1 vccd1 _1660_/X sky130_fd_sc_hd__and2_1
X_1591_ input76/X _1623_/A2 _1623_/B1 _2091_/Q hold521/X vssd1 vssd1 vccd1 vccd1 _1591_/X
+ sky130_fd_sc_hd__a221o_1
Xhold209 _1581_/X vssd1 vssd1 vccd1 vccd1 hold209/X sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_40_149 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__1167__A2 _1183_/A2 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_21_352 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_503 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_514 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_525 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_536 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_558 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_547 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_2212_ _2212_/CLK _2212_/D _1952_/Y vssd1 vssd1 vccd1 vccd1 _2212_/Q sky130_fd_sc_hd__dfrtp_4
XTAP_569 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_56_88 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_2143_ _2238_/CLK _2143_/D _1886_/Y vssd1 vssd1 vccd1 vccd1 _2143_/Q sky130_fd_sc_hd__dfrtp_2
X_2074_ _2106_/CLK _2074_/D _1817_/Y vssd1 vssd1 vccd1 vccd1 _2074_/Q sky130_fd_sc_hd__dfrtp_4
X_1025_ _1394_/B _1025_/B vssd1 vssd1 vccd1 vccd1 _1025_/Y sky130_fd_sc_hd__nor2_1
XFILLER_0_48_238 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_16_102 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_29_485 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_17_669 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_1927_ _1941_/A vssd1 vssd1 vccd1 vccd1 _1927_/Y sky130_fd_sc_hd__inv_2
XFILLER_0_44_477 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_4_530 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_21_80 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_1858_ _1949_/A vssd1 vssd1 vccd1 vccd1 _1858_/Y sky130_fd_sc_hd__inv_2
Xhold710 hold836/X vssd1 vssd1 vccd1 vccd1 hold710/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold721 hold860/X vssd1 vssd1 vccd1 vccd1 hold721/X sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_12_341 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xhold732 hold885/X vssd1 vssd1 vccd1 vccd1 hold732/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold743 hold743/A vssd1 vssd1 vccd1 vccd1 la_data_out[54] sky130_fd_sc_hd__buf_12
Xhold754 hold777/X vssd1 vssd1 vccd1 vccd1 hold754/X sky130_fd_sc_hd__dlygate4sd3_1
X_1789_ _2227_/Q _1802_/B vssd1 vssd1 vccd1 vccd1 _1789_/X sky130_fd_sc_hd__and2_1
XFILLER_0_40_650 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
Xhold776 _2145_/Q vssd1 vssd1 vccd1 vccd1 hold776/X sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA__1563__C1 hold136/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_12_374 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xhold765 _2158_/Q vssd1 vssd1 vccd1 vccd1 hold765/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold787 _2211_/Q vssd1 vssd1 vccd1 vccd1 hold787/X sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA_fanout583_A _1519_/B1 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xhold798 _2262_/Q vssd1 vssd1 vccd1 vccd1 hold798/X sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA__1094__A1 _2117_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_54_219 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_54_208 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_35_433 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_23_606 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_7_390 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__2062__A _2069_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_23_617 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_22_149 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XANTENNA__1149__A2 _1183_/A2 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_hold962_A _2098_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_30_193 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__1406__A _1415_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xhold70 hold70/A vssd1 vssd1 vccd1 vccd1 hold70/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold92 la_data_in[5] vssd1 vssd1 vccd1 vccd1 hold92/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold81 hold81/A vssd1 vssd1 vccd1 vccd1 hold81/X sky130_fd_sc_hd__buf_4
XFILLER_0_42_68 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_53_274 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_1712_ _2140_/Q _1802_/B vssd1 vssd1 vccd1 vccd1 _1712_/X sky130_fd_sc_hd__and2_1
XFILLER_0_5_349 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_26_477 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_1643_ _2071_/Q _1725_/B vssd1 vssd1 vccd1 vccd1 _1643_/X sky130_fd_sc_hd__and2_1
XANTENNA_1 _1400_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_1574_ hold291/X hold982/X hold81/X vssd1 vssd1 vccd1 vccd1 _2099_/D sky130_fd_sc_hd__mux2_1
XFILLER_0_21_160 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_311 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_300 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_322 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_333 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_344 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_355 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_366 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_388 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_377 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_399 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_2126_ _2223_/CLK _2126_/D _1869_/Y vssd1 vssd1 vccd1 vccd1 _2126_/Q sky130_fd_sc_hd__dfrtp_4
XPHY_17 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_2057_ _2069_/A vssd1 vssd1 vccd1 vccd1 _2057_/Y sky130_fd_sc_hd__inv_2
XPHY_28 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__1076__A1 _2126_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_1008_ _1198_/A _1811_/A vssd1 vssd1 vccd1 vccd1 _1008_/Y sky130_fd_sc_hd__nand2_1
XPHY_39 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_49_569 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_37_709 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_17_488 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_13_661 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_12_171 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xhold562 hold779/X vssd1 vssd1 vccd1 vccd1 _1191_/B sky130_fd_sc_hd__buf_1
Xhold540 hold540/A vssd1 vssd1 vccd1 vccd1 _0987_/B sky130_fd_sc_hd__dlygate4sd3_1
Xhold551 la_data_in[91] vssd1 vssd1 vccd1 vccd1 hold551/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold595 hold674/X vssd1 vssd1 vccd1 vccd1 hold595/X sky130_fd_sc_hd__dlymetal6s2s_1
Xhold584 hold688/X vssd1 vssd1 vccd1 vccd1 hold584/X sky130_fd_sc_hd__clkbuf_2
Xhold573 hold679/X vssd1 vssd1 vccd1 vccd1 hold573/X sky130_fd_sc_hd__clkbuf_2
XANTENNA__1551__A2 _1637_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__2057__A _2069_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__1067__B2 _1066_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__1896__A _2069_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_55_528 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_27_219 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_12_38 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_50_299 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_1290_ input39/X _1529_/A2 _1529_/B1 _2215_/Q hold285/X vssd1 vssd1 vccd1 vccd1 _1290_/X
+ sky130_fd_sc_hd__a221o_1
XFILLER_0_37_57 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xinput160 data_in[97] vssd1 vssd1 vccd1 vccd1 _1401_/A1 sky130_fd_sc_hd__buf_1
Xinput171 hold509/X vssd1 vssd1 vccd1 vccd1 hold510/A sky130_fd_sc_hd__buf_1
XFILLER_0_37_68 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
Xinput182 hold246/X vssd1 vssd1 vccd1 vccd1 hold247/A sky130_fd_sc_hd__clkbuf_1
Xinput193 hold342/X vssd1 vssd1 vccd1 vccd1 hold343/A sky130_fd_sc_hd__clkbuf_1
XFILLER_0_53_45 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_53_34 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_53_23 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_46_517 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_19_709 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_46_539 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_46_528 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_5_102 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_14_403 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__1230__A1 input61/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_14_469 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_1_330 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_1626_ hold177/X hold965/X _1632_/S vssd1 vssd1 vccd1 vccd1 _2073_/D sky130_fd_sc_hd__mux2_1
XFILLER_0_1_385 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_1557_ input94/X _1623_/A2 _1623_/B1 _2108_/Q hold336/X vssd1 vssd1 vccd1 vccd1 _1557_/X
+ sky130_fd_sc_hd__a221o_1
XTAP_130 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_141 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_1488_ hold349/X _2142_/Q _1504_/S vssd1 vssd1 vccd1 vccd1 _1488_/X sky130_fd_sc_hd__mux2_1
XTAP_174 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_152 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_163 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__1480__S _1504_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_196 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_185 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__1297__A1 _2212_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_2109_ _2177_/CLK _2109_/D _1852_/Y vssd1 vssd1 vccd1 vccd1 _2109_/Q sky130_fd_sc_hd__dfrtp_4
XANTENNA_fanout546_A _1792_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xclkbuf_1_0__f_wb_clk_i clkbuf_0_wb_clk_i/X vssd1 vssd1 vccd1 vccd1 clkbuf_leaf_9_wb_clk_i/A
+ sky130_fd_sc_hd__clkbuf_16
XFILLER_0_49_377 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_37_517 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_37_539 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_45_561 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_17_274 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_33_701 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_17_296 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XANTENNA_clkbuf_leaf_5_wb_clk_i_A clkbuf_leaf_9_wb_clk_i/A vssd1 vssd1 vccd1 vccd1
+ sky130_fd_sc_hd__diode_2
XANTENNA__1221__A1 input64/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xhold370 _1561_/X vssd1 vssd1 vccd1 vccd1 hold370/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold381 _1498_/X vssd1 vssd1 vccd1 vccd1 _2137_/D sky130_fd_sc_hd__dlygate4sd3_1
Xhold392 _1521_/X vssd1 vssd1 vccd1 vccd1 hold392/X sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA__1390__S _1435_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_hold925_A _2184_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__1288__A1 _2215_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_23_37 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_28_528 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xclkbuf_leaf_11_wb_clk_i clkbuf_1_1__f_wb_clk_i/X vssd1 vssd1 vccd1 vccd1 _2223_/CLK
+ sky130_fd_sc_hd__clkbuf_16
XANTENNA__1460__A1 _1527_/A2 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_24_701 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_36_583 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_36_594 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA_output465_A hold570/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_23_266 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__1212__A1 input68/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_23_277 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_1411_ _1410_/X _2174_/Q hold27/X vssd1 vssd1 vccd1 vccd1 _1411_/X sky130_fd_sc_hd__mux2_1
XANTENNA__1515__A2 _1519_/A2 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_1342_ _1341_/X _2197_/Q _1372_/S vssd1 vssd1 vccd1 vccd1 _1342_/X sky130_fd_sc_hd__mux2_1
X_1273_ _1272_/X _2220_/Q _1318_/S vssd1 vssd1 vccd1 vccd1 _1273_/X sky130_fd_sc_hd__mux2_1
XFILLER_0_59_620 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_59_642 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_42_531 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_14_222 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_0988_ _1012_/D _1012_/C vssd1 vssd1 vccd1 vccd1 _1014_/C sky130_fd_sc_hd__and2_2
XFILLER_0_30_704 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xoutput420 _1737_/X vssd1 vssd1 vccd1 vccd1 data_out[95] sky130_fd_sc_hd__buf_12
XFILLER_0_42_597 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_42_575 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_14_277 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
Xoutput442 hold766/X vssd1 vssd1 vccd1 vccd1 hold745/A sky130_fd_sc_hd__buf_6
Xoutput431 hold650/X vssd1 vssd1 vccd1 vccd1 la_data_out[104] sky130_fd_sc_hd__buf_12
Xoutput453 hold658/X vssd1 vssd1 vccd1 vccd1 la_data_out[38] sky130_fd_sc_hd__buf_12
Xoutput486 hold585/X vssd1 vssd1 vccd1 vccd1 la_data_out[71] sky130_fd_sc_hd__buf_12
Xoutput464 hold607/X vssd1 vssd1 vccd1 vccd1 la_data_out[49] sky130_fd_sc_hd__buf_12
Xoutput475 hold568/X vssd1 vssd1 vccd1 vccd1 la_data_out[60] sky130_fd_sc_hd__buf_12
X_1609_ input23/X _1637_/B _1635_/C _2082_/Q hold156/X vssd1 vssd1 vccd1 vccd1 _1609_/X
+ sky130_fd_sc_hd__a221o_1
Xoutput497 hold580/X vssd1 vssd1 vccd1 vccd1 la_data_out[82] sky130_fd_sc_hd__buf_12
XFILLER_0_49_163 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_45_391 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_18_583 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__1130__A0 _2191_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_55_122 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_1960_ _2002_/A vssd1 vssd1 vccd1 vccd1 _1960_/Y sky130_fd_sc_hd__inv_2
XFILLER_0_28_347 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_55_155 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_1891_ _1982_/A vssd1 vssd1 vccd1 vccd1 _1891_/Y sky130_fd_sc_hd__inv_2
XFILLER_0_43_328 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_24_531 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_59_11 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_11_214 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_24_575 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_11_258 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_1325_ _1349_/A _1325_/B vssd1 vssd1 vccd1 vccd1 _1325_/X sky130_fd_sc_hd__and2_1
X_1256_ _1277_/A _1256_/B vssd1 vssd1 vccd1 vccd1 _1256_/X sky130_fd_sc_hd__and2_1
XANTENNA__1121__B1 _1189_/B1 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_1187_ hold655/X _1189_/A2 _1189_/B1 _1186_/X vssd1 vssd1 vccd1 vccd1 _2251_/D sky130_fd_sc_hd__a22o_1
XFILLER_0_46_100 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_46_188 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_6_285 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_15_564 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_30_512 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_30_589 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
Xoutput283 _1760_/X vssd1 vssd1 vccd1 vccd1 data_out[118] sky130_fd_sc_hd__buf_12
Xoutput272 _1750_/X vssd1 vssd1 vccd1 vccd1 data_out[108] sky130_fd_sc_hd__buf_12
Xoutput294 _1770_/X vssd1 vssd1 vccd1 vccd1 data_out[128] sky130_fd_sc_hd__buf_12
XANTENNA__1112__A0 _2200_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__2065__A _2065_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_37_122 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_53_615 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_38_667 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_38_689 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA_hold992_A _2173_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_52_136 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_40_309 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__1179__B1 _1189_/B1 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__1409__A _1415_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_707 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_718 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_729 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_29_69 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_1110_ _2201_/Q _2109_/Q _1112_/S vssd1 vssd1 vccd1 vccd1 _1110_/X sky130_fd_sc_hd__mux2_1
X_2090_ _2182_/CLK _2090_/D _1833_/Y vssd1 vssd1 vccd1 vccd1 _2090_/Q sky130_fd_sc_hd__dfrtp_4
XFILLER_0_45_35 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_45_57 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_1041_ hold602/X _1057_/A2 _1057_/B1 _1040_/X vssd1 vssd1 vccd1 vccd1 _2324_/D sky130_fd_sc_hd__a22o_1
XFILLER_0_44_604 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_1943_ _1949_/A vssd1 vssd1 vccd1 vccd1 _1943_/Y sky130_fd_sc_hd__inv_2
XFILLER_0_28_155 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_44_648 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_43_125 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_1874_ _2002_/A vssd1 vssd1 vccd1 vccd1 _1874_/Y sky130_fd_sc_hd__inv_2
XFILLER_0_43_169 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
Xhold903 _2293_/Q vssd1 vssd1 vccd1 vccd1 hold903/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold925 _2184_/Q vssd1 vssd1 vccd1 vccd1 hold925/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold914 _2131_/Q vssd1 vssd1 vccd1 vccd1 hold914/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold936 _1345_/X vssd1 vssd1 vccd1 vccd1 _2196_/D sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_24_394 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
Xhold947 _2190_/Q vssd1 vssd1 vccd1 vccd1 hold947/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold969 _2095_/Q vssd1 vssd1 vccd1 vccd1 hold969/X sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_3_288 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
Xhold958 _2075_/Q vssd1 vssd1 vccd1 vccd1 hold958/X sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_36_3 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_1308_ input32/X _1197_/D _1541_/B1 _2209_/Q hold59/X vssd1 vssd1 vccd1 vccd1 hold60/A
+ sky130_fd_sc_hd__a221o_1
X_2288_ _2296_/CLK _2288_/D _2027_/Y vssd1 vssd1 vccd1 vccd1 _2288_/Q sky130_fd_sc_hd__dfrtp_1
X_1239_ input58/X _1495_/A2 _1495_/B1 _2232_/Q hold436/X vssd1 vssd1 vccd1 vccd1 _1239_/X
+ sky130_fd_sc_hd__a221o_1
XFILLER_0_47_475 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_47_453 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_47_442 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_19_155 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_22_309 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XANTENNA__1581__B1 _1623_/B1 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_30_397 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XANTENNA__1899__A _1949_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_15_49 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_53_401 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_38_475 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_41_629 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_1590_ hold530/X hold973/X hold81/X vssd1 vssd1 vccd1 vccd1 _2091_/D sky130_fd_sc_hd__mux2_1
XFILLER_0_21_386 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_504 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_515 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_526 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_537 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_548 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_2211_ _2256_/CLK _2211_/D _1951_/Y vssd1 vssd1 vccd1 vccd1 _2211_/Q sky130_fd_sc_hd__dfrtp_2
XTAP_559 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_2142_ _2224_/CLK _2142_/D _1885_/Y vssd1 vssd1 vccd1 vccd1 _2142_/Q sky130_fd_sc_hd__dfrtp_1
X_2073_ _2164_/CLK _2073_/D _1816_/Y vssd1 vssd1 vccd1 vccd1 _2073_/Q sky130_fd_sc_hd__dfrtp_4
X_1024_ _1385_/B _1382_/B _1376_/B _1379_/B vssd1 vssd1 vccd1 vccd1 _1198_/B sky130_fd_sc_hd__nor4_1
XANTENNA__1627__B2 _2073_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_17_637 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_16_136 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_1926_ _1941_/A vssd1 vssd1 vccd1 vccd1 _1926_/Y sky130_fd_sc_hd__inv_2
XFILLER_0_44_489 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_1857_ _1913_/A vssd1 vssd1 vccd1 vccd1 _1857_/Y sky130_fd_sc_hd__inv_2
Xhold700 hold806/X vssd1 vssd1 vccd1 vccd1 hold700/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold711 hold819/X vssd1 vssd1 vccd1 vccd1 hold711/X sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_31_128 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_1788_ _2226_/Q _1802_/B vssd1 vssd1 vccd1 vccd1 _1788_/X sky130_fd_sc_hd__and2_1
Xhold744 hold765/X vssd1 vssd1 vccd1 vccd1 hold766/A sky130_fd_sc_hd__buf_1
Xhold733 hold859/X vssd1 vssd1 vccd1 vccd1 hold733/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold755 _0969_/C vssd1 vssd1 vccd1 vccd1 hold755/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold722 hold824/X vssd1 vssd1 vccd1 vccd1 hold722/X sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA__1563__B1 _1569_/B1 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xhold766 hold766/A vssd1 vssd1 vccd1 vccd1 hold766/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold777 la_data_in[85] vssd1 vssd1 vccd1 vccd1 hold777/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold788 _2149_/Q vssd1 vssd1 vccd1 vccd1 hold788/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold799 _2258_/Q vssd1 vssd1 vccd1 vccd1 hold799/X sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA_fanout576_A _1201_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__1618__A1 _2077_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_50_415 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_23_629 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_31_673 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__1393__S _1435_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_hold955_A _2183_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_26_15 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
Xhold82 hold82/A vssd1 vssd1 vccd1 vccd1 hold82/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold71 hold71/A vssd1 vssd1 vccd1 vccd1 hold71/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold60 hold60/A vssd1 vssd1 vccd1 vccd1 hold60/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold93 hold93/A vssd1 vssd1 vccd1 vccd1 hold93/X sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA__1609__B2 _2082_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__1085__A2 _1095_/A2 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_42_47 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_38_272 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_53_242 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_1711_ _2139_/Q _1804_/B vssd1 vssd1 vccd1 vccd1 _1711_/X sky130_fd_sc_hd__and2_2
XFILLER_0_41_426 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA_2 la_data_in[21] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_1642_ _2070_/Q _1725_/B vssd1 vssd1 vccd1 vccd1 _1642_/X sky130_fd_sc_hd__and2_2
X_1573_ input85/X _1619_/A2 _1619_/B1 _2100_/Q hold290/X vssd1 vssd1 vccd1 vccd1 _1573_/X
+ sky130_fd_sc_hd__a221o_1
XANTENNA__1545__B1 _1545_/B1 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_22_673 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_312 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_301 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_323 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_334 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_345 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_356 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_367 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_389 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_378 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_2125_ _2217_/CLK _2125_/D _1868_/Y vssd1 vssd1 vccd1 vccd1 _2125_/Q sky130_fd_sc_hd__dfrtp_2
XPHY_18 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_2056_ _2069_/A vssd1 vssd1 vccd1 vccd1 _2056_/Y sky130_fd_sc_hd__inv_2
XPHY_29 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_49_559 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_1007_ _1007_/A _1007_/B vssd1 vssd1 vccd1 vccd1 _1811_/A sky130_fd_sc_hd__nand2_2
XANTENNA__1481__C1 hold515/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__1478__S _1504_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_29_294 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_1909_ _1922_/A vssd1 vssd1 vccd1 vccd1 _1909_/Y sky130_fd_sc_hd__inv_2
XFILLER_0_44_253 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_17_478 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_32_404 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_44_297 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xhold530 _1589_/X vssd1 vssd1 vccd1 vccd1 hold530/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold563 _1021_/X vssd1 vssd1 vccd1 vccd1 hold563/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold552 hold552/A vssd1 vssd1 vccd1 vccd1 _0992_/A sky130_fd_sc_hd__buf_1
Xhold541 _0973_/C vssd1 vssd1 vccd1 vccd1 _0971_/C sky130_fd_sc_hd__buf_2
Xhold596 hold685/X vssd1 vssd1 vccd1 vccd1 hold596/X sky130_fd_sc_hd__dlymetal6s2s_1
Xhold585 hold730/X vssd1 vssd1 vccd1 vccd1 hold585/X sky130_fd_sc_hd__dlymetal6s2s_1
Xhold574 hold681/X vssd1 vssd1 vccd1 vccd1 hold574/X sky130_fd_sc_hd__clkbuf_2
XTAP_890 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__1067__A2 _1095_/A2 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_27_209 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_36_710 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_35_231 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_51_713 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__1224__C1 hold443/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_35_297 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_50_256 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__1527__B1 _1527_/B1 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_31_492 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
Xinput161 data_in[98] vssd1 vssd1 vccd1 vccd1 _1398_/A1 sky130_fd_sc_hd__buf_1
Xinput150 data_in[88] vssd1 vssd1 vccd1 vccd1 _1428_/A1 sky130_fd_sc_hd__buf_1
Xinput172 hold508/X vssd1 vssd1 vccd1 vccd1 _1810_/A sky130_fd_sc_hd__buf_1
Xinput183 hold263/X vssd1 vssd1 vccd1 vccd1 hold236/A sky130_fd_sc_hd__clkbuf_1
Xinput194 hold334/X vssd1 vssd1 vccd1 vccd1 hold335/A sky130_fd_sc_hd__clkbuf_1
XFILLER_0_53_57 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_26_253 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_26_264 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__1215__C1 hold298/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_41_212 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_26_275 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_26_297 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__1230__A2 _1503_/A2 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_41_278 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_1_342 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_1625_ input97/X _1637_/B _1635_/C _2074_/Q hold176/X vssd1 vssd1 vccd1 vccd1 _1625_/X
+ sky130_fd_sc_hd__a221o_1
X_1556_ _1555_/X hold793/X hold80/X vssd1 vssd1 vccd1 vccd1 _2108_/D sky130_fd_sc_hd__mux2_1
XTAP_120 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_131 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_1487_ _1487_/A1 _1503_/A2 _1503_/B1 _2143_/Q hold348/X vssd1 vssd1 vccd1 vccd1 _1487_/X
+ sky130_fd_sc_hd__a221o_1
XTAP_175 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_153 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_142 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_164 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_197 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_186 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_2108_ _2177_/CLK _2108_/D _1851_/Y vssd1 vssd1 vccd1 vccd1 _2108_/Q sky130_fd_sc_hd__dfrtp_4
XFILLER_0_49_334 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA_fanout539_A hold79/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__1049__A2 _1095_/A2 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_2039_ _2039_/A vssd1 vssd1 vccd1 vccd1 _2039_/Y sky130_fd_sc_hd__inv_2
XFILLER_0_33_713 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_45_595 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__1221__A2 _1503_/A2 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_32_256 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__1509__B1 _1519_/B1 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xhold371 hold497/X vssd1 vssd1 vccd1 vccd1 hold371/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold360 _1242_/X vssd1 vssd1 vccd1 vccd1 hold360/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold393 _1522_/X vssd1 vssd1 vccd1 vccd1 _2125_/D sky130_fd_sc_hd__dlygate4sd3_1
Xhold382 hold397/X vssd1 vssd1 vccd1 vccd1 hold382/X sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA__2068__A _2069_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_55_304 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_23_49 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_24_713 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_23_223 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_1410_ _1410_/A1 _1569_/A2 _1201_/X _2175_/Q hold203/X vssd1 vssd1 vccd1 vccd1 _1410_/X
+ sky130_fd_sc_hd__a221o_1
X_1341_ input20/X _1533_/A2 _1533_/B1 _2198_/Q hold369/X vssd1 vssd1 vccd1 vccd1 _1341_/X
+ sky130_fd_sc_hd__a221o_1
X_1272_ input46/X _1519_/A2 _1519_/B1 _2221_/Q hold470/X vssd1 vssd1 vccd1 vccd1 _1272_/X
+ sky130_fd_sc_hd__a221o_1
XFILLER_0_59_698 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_58_164 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA_hold95_A hold95/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_58_197 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_6_401 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_54_370 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_0987_ _1453_/A _0987_/B _1453_/B _0987_/D vssd1 vssd1 vccd1 vccd1 _1012_/C sky130_fd_sc_hd__and4_1
Xoutput410 _1728_/X vssd1 vssd1 vccd1 vccd1 data_out[86] sky130_fd_sc_hd__buf_12
XFILLER_0_42_587 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_14_289 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
Xoutput421 _1738_/X vssd1 vssd1 vccd1 vccd1 data_out[96] sky130_fd_sc_hd__buf_12
Xoutput443 hold772/X vssd1 vssd1 vccd1 vccd1 hold753/A sky130_fd_sc_hd__buf_6
Xoutput432 hold596/X vssd1 vssd1 vccd1 vccd1 la_data_out[105] sky130_fd_sc_hd__buf_12
X_1608_ hold204/X hold932/X _1632_/S vssd1 vssd1 vccd1 vccd1 _2082_/D sky130_fd_sc_hd__mux2_1
Xoutput476 hold598/X vssd1 vssd1 vccd1 vccd1 la_data_out[61] sky130_fd_sc_hd__buf_12
Xoutput487 hold621/X vssd1 vssd1 vccd1 vccd1 la_data_out[72] sky130_fd_sc_hd__buf_12
Xoutput454 hold623/X vssd1 vssd1 vccd1 vccd1 la_data_out[39] sky130_fd_sc_hd__buf_12
Xoutput465 hold570/X vssd1 vssd1 vccd1 vccd1 la_data_out[50] sky130_fd_sc_hd__buf_12
Xoutput498 hold653/X vssd1 vssd1 vccd1 vccd1 la_data_out[83] sky130_fd_sc_hd__buf_12
X_1539_ _1539_/A1 _1197_/D _1541_/B1 _2117_/Q hold59/X vssd1 vssd1 vccd1 vccd1 _1539_/X
+ sky130_fd_sc_hd__a221o_1
XFILLER_0_37_304 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_52_307 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_18_540 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_20_204 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xhold190 hold190/A vssd1 vssd1 vccd1 vccd1 _1325_/B sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_18_16 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__1130__A1 _2099_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_34_15 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_34_37 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_1890_ _1979_/A vssd1 vssd1 vccd1 vccd1 _1890_/Y sky130_fd_sc_hd__inv_2
XFILLER_0_3_415 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_51_373 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_24_587 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_51_384 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_1324_ _1323_/X _2203_/Q hold27/X vssd1 vssd1 vccd1 vccd1 _1324_/X sky130_fd_sc_hd__mux2_1
X_1255_ hold318/X hold904/X hold26/X vssd1 vssd1 vccd1 vccd1 _2226_/D sky130_fd_sc_hd__mux2_1
XANTENNA__1121__B2 _1120_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_1186_ _2163_/Q _2071_/Q _1188_/S vssd1 vssd1 vccd1 vccd1 _1186_/X sky130_fd_sc_hd__mux2_1
XFILLER_0_19_326 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_19_337 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_46_145 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_27_381 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__1486__S _1504_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_42_340 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__1188__A1 _2070_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_30_502 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_30_557 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xoutput273 _1751_/X vssd1 vssd1 vccd1 vccd1 data_out[109] sky130_fd_sc_hd__buf_12
Xoutput295 _1771_/X vssd1 vssd1 vccd1 vccd1 data_out[129] sky130_fd_sc_hd__buf_12
Xoutput284 _1761_/X vssd1 vssd1 vccd1 vccd1 data_out[119] sky130_fd_sc_hd__buf_12
XANTENNA__1360__A1 _2191_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__1112__A1 _2108_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_52_115 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__1396__S _1435_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_37_178 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA_hold985_A _2087_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_29_15 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_719 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_708 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_1040_ _2236_/Q _2144_/Q _1094_/S vssd1 vssd1 vccd1 vccd1 _1040_/X sky130_fd_sc_hd__mux2_1
XFILLER_0_29_613 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_1942_ _1949_/A vssd1 vssd1 vccd1 vccd1 _1942_/Y sky130_fd_sc_hd__inv_2
XFILLER_0_29_668 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_29_679 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_1873_ _2002_/A vssd1 vssd1 vccd1 vccd1 _1873_/Y sky130_fd_sc_hd__inv_2
XFILLER_0_44_638 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_43_137 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_4_713 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xhold904 _2226_/Q vssd1 vssd1 vccd1 vccd1 hold904/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold937 _2101_/Q vssd1 vssd1 vccd1 vccd1 hold937/X sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_51_181 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
Xhold926 _2189_/Q vssd1 vssd1 vccd1 vccd1 hold926/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold915 la_data_in[29] vssd1 vssd1 vccd1 vccd1 hold915/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold959 _2194_/Q vssd1 vssd1 vccd1 vccd1 hold959/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold948 _2200_/Q vssd1 vssd1 vccd1 vccd1 hold948/X sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA__1342__A1 _2197_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_1307_ _1310_/A hold58/X vssd1 vssd1 vccd1 vccd1 hold59/A sky130_fd_sc_hd__and2_1
X_2287_ _2300_/CLK _2287_/D _2026_/Y vssd1 vssd1 vccd1 vccd1 _2287_/Q sky130_fd_sc_hd__dfrtp_1
X_1238_ _1271_/A _1238_/B vssd1 vssd1 vccd1 vccd1 _1238_/X sky130_fd_sc_hd__and2_1
XFILLER_0_29_3 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_1169_ hold627/X _1183_/A2 _1183_/B1 _1168_/X vssd1 vssd1 vccd1 vccd1 _2260_/D sky130_fd_sc_hd__a22o_1
XFILLER_0_59_281 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA_fanout521_A hold26/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_35_605 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_19_167 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_34_137 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_30_354 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__1581__B2 _2096_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__1097__B1 _1097_/B1 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_38_421 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_26_616 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_505 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_516 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_2210_ _2212_/CLK _2210_/D _1950_/Y vssd1 vssd1 vccd1 vccd1 _2210_/Q sky130_fd_sc_hd__dfrtp_4
XTAP_527 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_538 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_549 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_56_46 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__1324__A1 _2203_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_2141_ _2238_/CLK _2141_/D _1884_/Y vssd1 vssd1 vccd1 vccd1 _2141_/Q sky130_fd_sc_hd__dfrtp_1
X_2072_ _2164_/CLK hold19/X _1815_/Y vssd1 vssd1 vccd1 vccd1 _2072_/Q sky130_fd_sc_hd__dfrtp_4
X_1023_ _1805_/A _1811_/A vssd1 vssd1 vccd1 vccd1 _1023_/Y sky130_fd_sc_hd__nor2_2
XANTENNA__1088__A0 _2212_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__1627__A2 _1637_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_29_443 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_56_251 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xclkbuf_leaf_6_wb_clk_i clkbuf_leaf_9_wb_clk_i/A vssd1 vssd1 vccd1 vccd1 _2194_/CLK
+ sky130_fd_sc_hd__clkbuf_16
X_1925_ _1941_/A vssd1 vssd1 vccd1 vccd1 _1925_/Y sky130_fd_sc_hd__inv_2
XFILLER_0_44_435 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__1260__B1 _1519_/B1 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_44_468 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_1856_ _1913_/A vssd1 vssd1 vccd1 vccd1 _1856_/Y sky130_fd_sc_hd__inv_2
XFILLER_0_25_671 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_1787_ _2225_/Q _1798_/B vssd1 vssd1 vccd1 vccd1 _1787_/X sky130_fd_sc_hd__and2_1
Xhold701 hold837/X vssd1 vssd1 vccd1 vccd1 hold701/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold712 hold826/X vssd1 vssd1 vccd1 vccd1 hold712/X sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_25_682 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
Xhold745 hold745/A vssd1 vssd1 vccd1 vccd1 la_data_out[123] sky130_fd_sc_hd__buf_12
XFILLER_0_4_587 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xhold734 hold868/X vssd1 vssd1 vccd1 vccd1 hold734/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold723 hold830/X vssd1 vssd1 vccd1 vccd1 hold723/X sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_24_192 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_40_641 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__1563__B2 _2105_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_12_387 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
Xhold756 _1451_/X vssd1 vssd1 vccd1 vccd1 hold90/A sky130_fd_sc_hd__dlygate4sd3_1
Xhold767 _2157_/Q vssd1 vssd1 vccd1 vccd1 hold767/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold778 _1018_/Y vssd1 vssd1 vccd1 vccd1 hold778/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold789 _1030_/X vssd1 vssd1 vccd1 vccd1 hold789/X sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA__1079__B1 _1095_/B1 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_39_207 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_35_402 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_16_660 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_22_129 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_15_192 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_31_641 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XANTENNA__1306__A1 _2209_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_hold948_A _2200_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xhold50 hold50/A vssd1 vssd1 vccd1 vccd1 hold50/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold83 hold98/X vssd1 vssd1 vccd1 vccd1 hold83/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold72 hold72/A vssd1 vssd1 vccd1 vccd1 hold72/X sky130_fd_sc_hd__buf_1
XFILLER_0_26_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xhold61 hold61/A vssd1 vssd1 vccd1 vccd1 hold61/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold94 hold94/A vssd1 vssd1 vccd1 vccd1 hold94/X sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA__1609__A2 _1637_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_42_15 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_5_318 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_38_284 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_38_295 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_53_254 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_14_619 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_1710_ _2138_/Q _1804_/B vssd1 vssd1 vccd1 vccd1 _1710_/X sky130_fd_sc_hd__and2_2
XFILLER_0_41_449 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_1641_ _2157_/Q _1810_/C vssd1 vssd1 vccd1 vccd1 _1641_/Y sky130_fd_sc_hd__nor2_1
XANTENNA_3 la_data_in[22] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_22_641 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_1572_ _1571_/X hold929/X hold81/X vssd1 vssd1 vccd1 vccd1 _2100_/D sky130_fd_sc_hd__mux2_1
XANTENNA__1545__B2 _2114_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_21_151 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_313 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_302 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_324 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_335 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_346 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_357 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_368 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_379 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_2124_ _2217_/CLK _2124_/D _1867_/Y vssd1 vssd1 vccd1 vccd1 _2124_/Q sky130_fd_sc_hd__dfrtp_2
XFILLER_0_49_505 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_2055_ _2069_/A vssd1 vssd1 vccd1 vccd1 _2055_/Y sky130_fd_sc_hd__inv_2
XPHY_19 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_1006_ _1367_/B _1364_/B _1370_/B _1373_/B vssd1 vssd1 vccd1 vccd1 _1007_/B sky130_fd_sc_hd__and4b_1
XFILLER_0_16_82 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__1481__B1 _1503_/B1 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_29_240 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__1233__B1 _1503_/B1 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_44_265 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_1908_ _1922_/A vssd1 vssd1 vccd1 vccd1 _1908_/Y sky130_fd_sc_hd__inv_2
XFILLER_0_17_457 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_1839_ _1922_/A vssd1 vssd1 vccd1 vccd1 _1839_/Y sky130_fd_sc_hd__inv_2
XFILLER_0_4_340 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
Xhold520 _1808_/C vssd1 vssd1 vccd1 vccd1 _1385_/B sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA__1494__S _1504_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xhold553 _1012_/B vssd1 vssd1 vccd1 vccd1 _0993_/D sky130_fd_sc_hd__dlygate4sd3_1
Xhold542 _0975_/Y vssd1 vssd1 vccd1 vccd1 _0986_/A sky130_fd_sc_hd__buf_1
Xhold531 la_data_in[20] vssd1 vssd1 vccd1 vccd1 hold531/X sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA__1536__A1 _2118_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xhold564 _1022_/B vssd1 vssd1 vccd1 vccd1 _1466_/S sky130_fd_sc_hd__clkbuf_2
Xhold597 hold719/X vssd1 vssd1 vccd1 vccd1 hold597/X sky130_fd_sc_hd__dlymetal6s2s_1
Xhold586 hold701/X vssd1 vssd1 vccd1 vccd1 hold586/X sky130_fd_sc_hd__clkbuf_2
Xhold575 hold666/X vssd1 vssd1 vccd1 vccd1 hold575/X sky130_fd_sc_hd__dlymetal6s2s_1
XTAP_880 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_891 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__1472__A0 _1471_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__1224__B1 _1503_/B1 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xcontroller_650 vssd1 vssd1 vccd1 vccd1 controller_650/HI la_data_out[114] sky130_fd_sc_hd__conb_1
XFILLER_0_23_427 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_50_246 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_23_449 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_50_279 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XANTENNA__1527__B2 _2123_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__1527__A1 _1527_/A1 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_37_15 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
Xinput162 data_in[99] vssd1 vssd1 vccd1 vccd1 _1395_/A1 sky130_fd_sc_hd__clkbuf_1
Xinput140 data_in[79] vssd1 vssd1 vccd1 vccd1 _1473_/A1 sky130_fd_sc_hd__buf_2
Xinput151 data_in[89] vssd1 vssd1 vccd1 vccd1 _1425_/A1 sky130_fd_sc_hd__clkbuf_1
Xinput173 hold504/X vssd1 vssd1 vccd1 vccd1 hold88/A sky130_fd_sc_hd__buf_1
Xinput184 hold221/X vssd1 vssd1 vccd1 vccd1 hold222/A sky130_fd_sc_hd__clkbuf_1
Xinput195 hold225/X vssd1 vssd1 vccd1 vccd1 hold226/A sky130_fd_sc_hd__clkbuf_1
XFILLER_0_53_69 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_27_711 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_26_232 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_1624_ _1623_/X hold951/X _1632_/S vssd1 vssd1 vccd1 vccd1 _1624_/X sky130_fd_sc_hd__mux2_1
XFILLER_0_1_354 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_1555_ input95/X _1637_/B _1635_/C _2109_/Q hold227/X vssd1 vssd1 vccd1 vccd1 _1555_/X
+ sky130_fd_sc_hd__a221o_1
XTAP_121 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_132 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_1486_ hold423/X hold910/X _1504_/S vssd1 vssd1 vccd1 vccd1 _2143_/D sky130_fd_sc_hd__mux2_1
XFILLER_0_10_699 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_154 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_143 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_165 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_198 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_187 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_176 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__1343__A _1415_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_2107_ _2177_/CLK _2107_/D _1850_/Y vssd1 vssd1 vccd1 vccd1 _2107_/Q sky130_fd_sc_hd__dfrtp_4
XFILLER_0_11_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_2038_ _2061_/A vssd1 vssd1 vccd1 vccd1 _2038_/Y sky130_fd_sc_hd__inv_2
XFILLER_0_45_574 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_17_265 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA_fanout601_A _1922_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_17_287 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__1509__A1 _1509_/A1 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_20_408 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
Xhold350 _1488_/X vssd1 vssd1 vccd1 vccd1 _2142_/D sky130_fd_sc_hd__dlygate4sd3_1
Xhold361 _1243_/X vssd1 vssd1 vccd1 vccd1 _2230_/D sky130_fd_sc_hd__dlygate4sd3_1
Xhold383 hold383/A vssd1 vssd1 vccd1 vccd1 _1232_/B sky130_fd_sc_hd__dlygate4sd3_1
Xhold372 hold372/A vssd1 vssd1 vccd1 vccd1 _1262_/B sky130_fd_sc_hd__dlygate4sd3_1
Xhold394 hold883/X vssd1 vssd1 vccd1 vccd1 hold394/X sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA__1700__B _1715_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__1399__S _1435_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_36_530 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_11_419 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_1340_ _1349_/A _1340_/B vssd1 vssd1 vccd1 vccd1 _1340_/X sky130_fd_sc_hd__and2_1
XFILLER_0_31_290 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xclkbuf_leaf_20_wb_clk_i clkbuf_1_1__f_wb_clk_i/X vssd1 vssd1 vccd1 vccd1 _2328_/CLK
+ sky130_fd_sc_hd__clkbuf_16
X_1271_ _1271_/A _1271_/B vssd1 vssd1 vccd1 vccd1 _1271_/X sky130_fd_sc_hd__and2_1
XANTENNA__1102__S _1112_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_19_519 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_54_382 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_42_511 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_0986_ _0986_/A _0986_/B vssd1 vssd1 vccd1 vccd1 _0986_/Y sky130_fd_sc_hd__nor2_1
XFILLER_0_42_544 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_42_533 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
Xoutput411 _1729_/X vssd1 vssd1 vccd1 vccd1 data_out[87] sky130_fd_sc_hd__buf_12
Xoutput400 _1719_/X vssd1 vssd1 vccd1 vccd1 data_out[77] sky130_fd_sc_hd__buf_12
Xoutput422 _1739_/X vssd1 vssd1 vccd1 vccd1 data_out[97] sky130_fd_sc_hd__buf_12
Xoutput444 hold770/X vssd1 vssd1 vccd1 vccd1 hold751/A sky130_fd_sc_hd__buf_6
Xoutput433 hold602/X vssd1 vssd1 vccd1 vccd1 la_data_out[106] sky130_fd_sc_hd__buf_12
X_1607_ input34/X _1623_/A2 _1623_/B1 _2083_/Q hold203/X vssd1 vssd1 vccd1 vccd1 _1607_/X
+ sky130_fd_sc_hd__a221o_1
XFILLER_0_59_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
Xoutput477 hold612/X vssd1 vssd1 vccd1 vccd1 la_data_out[62] sky130_fd_sc_hd__buf_12
Xoutput466 hold626/X vssd1 vssd1 vccd1 vccd1 la_data_out[51] sky130_fd_sc_hd__buf_12
Xoutput455 hold638/X vssd1 vssd1 vccd1 vccd1 la_data_out[40] sky130_fd_sc_hd__buf_12
Xoutput499 hold652/X vssd1 vssd1 vccd1 vccd1 la_data_out[84] sky130_fd_sc_hd__buf_12
Xoutput488 hold746/X vssd1 vssd1 vccd1 vccd1 hold747/A sky130_fd_sc_hd__buf_6
X_1538_ _1537_/X _2117_/Q hold80/X vssd1 vssd1 vccd1 vccd1 _1538_/X sky130_fd_sc_hd__mux2_1
X_1469_ _1469_/A1 _1197_/D hold7/X vssd1 vssd1 vccd1 vccd1 hold8/A sky130_fd_sc_hd__a21o_1
XANTENNA_fanout551_A _1641_/Y vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_18_596 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_33_500 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_45_393 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_33_544 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_20_249 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xhold180 hold881/X vssd1 vssd1 vccd1 vccd1 hold70/A sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_0_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xhold191 _1325_/X vssd1 vssd1 vccd1 vccd1 hold191/X sky130_fd_sc_hd__buf_1
XANTENNA_hold930_A _2119_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_50_15 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_36_360 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_3_405 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_24_533 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XANTENNA_clkbuf_leaf_19_wb_clk_i_A clkbuf_1_1__f_wb_clk_i/X vssd1 vssd1 vccd1 vccd1
+ sky130_fd_sc_hd__diode_2
XFILLER_0_59_57 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_11_238 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_1323_ input27/X _1197_/D _1541_/B1 _2204_/Q hold183/X vssd1 vssd1 vccd1 vccd1 _1323_/X
+ sky130_fd_sc_hd__a221o_1
X_1254_ input52/X _1503_/A2 _1503_/B1 _2227_/Q hold317/X vssd1 vssd1 vccd1 vccd1 _1254_/X
+ sky130_fd_sc_hd__a221o_1
XANTENNA__1121__A2 _1189_/A2 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_1185_ hold603/X _1189_/A2 _1189_/B1 _1184_/X vssd1 vssd1 vccd1 vccd1 _2252_/D sky130_fd_sc_hd__a22o_1
XFILLER_0_59_474 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_59_452 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_46_124 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_0969_ _0977_/D _0971_/C _0969_/C vssd1 vssd1 vccd1 vccd1 _1197_/A sky130_fd_sc_hd__nor3_1
XFILLER_0_27_393 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_40_81 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__1593__C1 _1388_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_30_547 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA_fanout599_A input262/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xoutput285 _1653_/X vssd1 vssd1 vccd1 vccd1 data_out[11] sky130_fd_sc_hd__buf_12
Xoutput263 _1642_/X vssd1 vssd1 vccd1 vccd1 data_out[0] sky130_fd_sc_hd__buf_12
Xoutput274 _1652_/X vssd1 vssd1 vccd1 vccd1 data_out[10] sky130_fd_sc_hd__buf_12
Xoutput296 _1654_/X vssd1 vssd1 vccd1 vccd1 data_out[12] sky130_fd_sc_hd__buf_12
XFILLER_0_38_658 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_33_330 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__1179__A2 _1189_/A2 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_hold978_A _2195_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_709 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_29_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_45_26 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_45_15 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_28_113 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_1941_ _1941_/A vssd1 vssd1 vccd1 vccd1 _1941_/Y sky130_fd_sc_hd__inv_2
X_1872_ _2002_/A vssd1 vssd1 vccd1 vccd1 _1872_/Y sky130_fd_sc_hd__inv_2
XFILLER_0_37_680 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_43_149 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_37_691 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xhold916 _1360_/X vssd1 vssd1 vccd1 vccd1 _2191_/D sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA__1575__C1 hold223/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xhold905 _2307_/Q vssd1 vssd1 vccd1 vccd1 hold905/X sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_24_374 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xhold927 _2094_/Q vssd1 vssd1 vccd1 vccd1 hold927/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold938 _2096_/Q vssd1 vssd1 vccd1 vccd1 hold938/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold949 _2176_/Q vssd1 vssd1 vccd1 vccd1 hold949/X sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_20_580 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_1306_ hold96/X _2209_/Q _1318_/S vssd1 vssd1 vccd1 vccd1 hold97/A sky130_fd_sc_hd__mux2_1
X_2286_ _2300_/CLK _2286_/D _2025_/Y vssd1 vssd1 vccd1 vccd1 _2286_/Q sky130_fd_sc_hd__dfrtp_1
X_1237_ _1236_/X _2232_/Q _1252_/S vssd1 vssd1 vccd1 vccd1 _1237_/X sky130_fd_sc_hd__mux2_1
X_1168_ hold988/X _2080_/Q _1188_/S vssd1 vssd1 vccd1 vccd1 _1168_/X sky130_fd_sc_hd__mux2_1
XFILLER_0_47_400 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_1099_ hold566/X _1157_/A2 _1157_/B1 _1098_/X vssd1 vssd1 vccd1 vccd1 _2295_/D sky130_fd_sc_hd__a22o_1
XFILLER_0_34_105 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_35_617 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_35_628 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_42_193 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__1581__A2 _1623_/A2 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_25_116 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_38_477 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_506 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_517 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_528 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_539 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_56_25 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_2140_ _2239_/CLK _2140_/D _1883_/Y vssd1 vssd1 vccd1 vccd1 _2140_/Q sky130_fd_sc_hd__dfrtp_1
X_2071_ _2164_/CLK hold33/X _1814_/Y vssd1 vssd1 vccd1 vccd1 _2071_/Q sky130_fd_sc_hd__dfrtp_4
X_1022_ _1277_/A _1022_/B vssd1 vssd1 vccd1 vccd1 _1022_/X sky130_fd_sc_hd__or2_1
XANTENNA__1088__A1 _2120_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_1924_ _1941_/A vssd1 vssd1 vccd1 vccd1 _1924_/Y sky130_fd_sc_hd__inv_2
XFILLER_0_8_338 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_17_617 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_29_466 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_29_477 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__1260__A1 input50/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_4_500 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_16_127 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__1110__S _1112_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_1855_ _1988_/A vssd1 vssd1 vccd1 vccd1 _1855_/Y sky130_fd_sc_hd__inv_2
X_1786_ _2224_/Q _1798_/B vssd1 vssd1 vccd1 vccd1 _1786_/X sky130_fd_sc_hd__and2_1
Xhold702 hold762/X vssd1 vssd1 vccd1 vccd1 hold702/X sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_21_83 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_25_694 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_40_631 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_12_344 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
Xhold724 hold833/X vssd1 vssd1 vccd1 vccd1 hold724/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold746 hold763/X vssd1 vssd1 vccd1 vccd1 hold746/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold735 hold838/X vssd1 vssd1 vccd1 vccd1 hold735/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold713 hold821/X vssd1 vssd1 vccd1 vccd1 hold713/X sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA__1563__A2 _1569_/A2 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xhold768 hold768/A vssd1 vssd1 vccd1 vccd1 hold768/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold757 _1452_/X vssd1 vssd1 vccd1 vccd1 hold91/A sky130_fd_sc_hd__dlygate4sd3_1
Xhold779 _1204_/B vssd1 vssd1 vccd1 vccd1 hold779/X sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA__1346__A _1415_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_41_3 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_2269_ _2269_/CLK _2269_/D _2008_/Y vssd1 vssd1 vccd1 vccd1 _2269_/Q sky130_fd_sc_hd__dfrtp_1
XANTENNA__1079__B2 _1078_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_39_219 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__1251__A1 input53/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_7_371 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_43_480 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_16_672 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_16_694 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_31_653 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_30_141 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
Xhold40 hold40/A vssd1 vssd1 vccd1 vccd1 hold40/X sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA__1703__B _1715_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xhold62 hold62/A vssd1 vssd1 vccd1 vccd1 hold62/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold51 hold51/A vssd1 vssd1 vccd1 vccd1 hold51/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold73 hold73/A vssd1 vssd1 vccd1 vccd1 hold73/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold84 hold84/A vssd1 vssd1 vccd1 vccd1 hold84/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold95 hold95/A vssd1 vssd1 vccd1 vccd1 hold95/X sky130_fd_sc_hd__buf_1
XFILLER_0_42_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_26_425 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__1242__A1 input57/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_53_299 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_1640_ _2156_/Q _1455_/A _1637_/B _0955_/Y _1635_/C vssd1 vssd1 vccd1 vccd1 _2249_/D
+ sky130_fd_sc_hd__a221o_1
XFILLER_0_34_480 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_1571_ input87/X _1623_/A2 _1623_/B1 _2101_/Q hold276/X vssd1 vssd1 vccd1 vccd1 _1571_/X
+ sky130_fd_sc_hd__a221o_1
XANTENNA_4 la_data_in[23] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_21_130 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_314 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_303 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_325 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_336 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_347 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_358 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_369 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_2123_ _2217_/CLK _2123_/D _1866_/Y vssd1 vssd1 vccd1 vccd1 _2123_/Q sky130_fd_sc_hd__dfrtp_2
X_2054_ _2061_/A vssd1 vssd1 vccd1 vccd1 _2054_/Y sky130_fd_sc_hd__inv_2
X_1005_ _1361_/B _1355_/B _1352_/B _1358_/B vssd1 vssd1 vccd1 vccd1 _1007_/A sky130_fd_sc_hd__and4bb_1
XANTENNA__1481__A1 _1481_/A1 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_57_561 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_8_179 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_32_82 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__1233__A1 input60/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_1907_ _1916_/A vssd1 vssd1 vccd1 vccd1 _1907_/Y sky130_fd_sc_hd__inv_2
XFILLER_0_4_352 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_1838_ _1852_/A vssd1 vssd1 vccd1 vccd1 _1838_/Y sky130_fd_sc_hd__inv_2
Xhold510 hold510/A vssd1 vssd1 vccd1 vccd1 _1025_/B sky130_fd_sc_hd__buf_1
Xhold554 _0993_/X vssd1 vssd1 vccd1 vccd1 hold554/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold543 _0986_/Y vssd1 vssd1 vccd1 vccd1 _1192_/C sky130_fd_sc_hd__buf_1
Xhold532 la_data_in[21] vssd1 vssd1 vccd1 vccd1 hold532/X sky130_fd_sc_hd__dlygate4sd3_1
X_1769_ _2207_/Q _1804_/B vssd1 vssd1 vccd1 vccd1 _1769_/X sky130_fd_sc_hd__and2_1
Xhold521 _1385_/X vssd1 vssd1 vccd1 vccd1 hold521/X sky130_fd_sc_hd__dlymetal6s2s_1
XFILLER_0_40_461 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xhold587 hold696/X vssd1 vssd1 vccd1 vccd1 hold587/X sky130_fd_sc_hd__buf_1
Xhold565 _1145_/X vssd1 vssd1 vccd1 vccd1 _2272_/D sky130_fd_sc_hd__dlygate4sd3_1
Xhold576 hold704/X vssd1 vssd1 vccd1 vccd1 hold576/X sky130_fd_sc_hd__clkbuf_2
Xhold598 hold708/X vssd1 vssd1 vccd1 vccd1 hold598/X sky130_fd_sc_hd__dlymetal6s2s_1
XTAP_870 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_892 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_881 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_36_701 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_35_222 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__1224__A1 input63/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xcontroller_651 vssd1 vssd1 vccd1 vccd1 controller_651/HI la_data_out[115] sky130_fd_sc_hd__conb_1
Xcontroller_640 vssd1 vssd1 vccd1 vccd1 controller_640/HI la_data_out[22] sky130_fd_sc_hd__conb_1
XFILLER_0_35_266 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_23_439 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA_hold793_A _2108_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__1527__A2 _1527_/A2 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_31_472 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_37_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
Xinput152 data_in[8] vssd1 vssd1 vccd1 vccd1 _1615_/A1 sky130_fd_sc_hd__buf_1
Xinput130 data_in[6] vssd1 vssd1 vccd1 vccd1 _1619_/A1 sky130_fd_sc_hd__clkbuf_1
Xinput163 data_in[9] vssd1 vssd1 vccd1 vccd1 _1613_/A1 sky130_fd_sc_hd__buf_1
Xinput141 data_in[7] vssd1 vssd1 vccd1 vccd1 _1617_/A1 sky130_fd_sc_hd__clkbuf_1
Xinput196 hold252/X vssd1 vssd1 vccd1 vccd1 hold253/A sky130_fd_sc_hd__clkbuf_1
Xinput174 hold458/X vssd1 vssd1 vccd1 vccd1 hold2/A sky130_fd_sc_hd__buf_1
Xinput185 hold288/X vssd1 vssd1 vccd1 vccd1 hold289/A sky130_fd_sc_hd__clkbuf_1
XANTENNA__1160__A0 _2176_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_53_15 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_53_48 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_39_561 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_26_222 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_26_244 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__1215__A1 input66/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_54_586 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_41_225 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_22_450 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_1623_ _1623_/A1 _1623_/A2 _1623_/B1 _2075_/Q hold281/X vssd1 vssd1 vccd1 vccd1 _1623_/X
+ sky130_fd_sc_hd__a221o_1
XFILLER_0_1_366 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_1554_ _1553_/X hold786/X _1632_/S vssd1 vssd1 vccd1 vccd1 _2109_/D sky130_fd_sc_hd__mux2_1
X_1485_ _1485_/A1 _1503_/A2 _1503_/B1 _2144_/Q hold422/X vssd1 vssd1 vccd1 vccd1 _1485_/X
+ sky130_fd_sc_hd__a221o_1
XTAP_122 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_133 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_155 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_144 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_166 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
.ends

