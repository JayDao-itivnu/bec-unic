VERSION 5.7 ;
  NOWIREEXTENSIONATPIN ON ;
  DIVIDERCHAR "/" ;
  BUSBITCHARS "[]" ;
MACRO sm_bec_v3
  CLASS BLOCK ;
  FOREIGN sm_bec_v3 ;
  ORIGIN 0.000 0.000 ;
  SIZE 579.150 BY 589.870 ;
  PIN becStatus[0]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 2.673000 ;
    PORT
      LAYER met3 ;
        RECT 0.000 511.400 4.000 512.000 ;
    END
  END becStatus[0]
  PIN becStatus[1]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 2.673000 ;
    PORT
      LAYER met3 ;
        RECT 0.000 514.120 4.000 514.720 ;
    END
  END becStatus[1]
  PIN becStatus[2]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 2.673000 ;
    PORT
      LAYER met3 ;
        RECT 0.000 516.840 4.000 517.440 ;
    END
  END becStatus[2]
  PIN becStatus[3]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 2.673000 ;
    PORT
      LAYER met3 ;
        RECT 0.000 519.560 4.000 520.160 ;
    END
  END becStatus[3]
  PIN clk
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.852000 ;
    ANTENNADIFFAREA 0.434700 ;
    PORT
      LAYER met2 ;
        RECT 48.850 0.000 49.130 4.000 ;
    END
  END clk
  PIN data_in[0]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.126000 ;
    ANTENNADIFFAREA 0.434700 ;
    PORT
      LAYER met3 ;
        RECT 575.150 69.400 579.150 70.000 ;
    END
  END data_in[0]
  PIN data_in[100]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.126000 ;
    ANTENNADIFFAREA 0.434700 ;
    PORT
      LAYER met3 ;
        RECT 575.150 341.400 579.150 342.000 ;
    END
  END data_in[100]
  PIN data_in[101]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.126000 ;
    ANTENNADIFFAREA 0.434700 ;
    PORT
      LAYER met3 ;
        RECT 575.150 344.120 579.150 344.720 ;
    END
  END data_in[101]
  PIN data_in[102]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.126000 ;
    ANTENNADIFFAREA 0.434700 ;
    PORT
      LAYER met3 ;
        RECT 575.150 346.840 579.150 347.440 ;
    END
  END data_in[102]
  PIN data_in[103]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.126000 ;
    ANTENNADIFFAREA 0.434700 ;
    PORT
      LAYER met3 ;
        RECT 575.150 349.560 579.150 350.160 ;
    END
  END data_in[103]
  PIN data_in[104]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.126000 ;
    ANTENNADIFFAREA 0.434700 ;
    PORT
      LAYER met3 ;
        RECT 575.150 352.280 579.150 352.880 ;
    END
  END data_in[104]
  PIN data_in[105]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.126000 ;
    ANTENNADIFFAREA 0.434700 ;
    PORT
      LAYER met3 ;
        RECT 575.150 355.000 579.150 355.600 ;
    END
  END data_in[105]
  PIN data_in[106]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.126000 ;
    ANTENNADIFFAREA 0.434700 ;
    PORT
      LAYER met3 ;
        RECT 575.150 357.720 579.150 358.320 ;
    END
  END data_in[106]
  PIN data_in[107]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.126000 ;
    ANTENNADIFFAREA 0.434700 ;
    PORT
      LAYER met3 ;
        RECT 575.150 360.440 579.150 361.040 ;
    END
  END data_in[107]
  PIN data_in[108]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.126000 ;
    ANTENNADIFFAREA 0.434700 ;
    PORT
      LAYER met3 ;
        RECT 575.150 363.160 579.150 363.760 ;
    END
  END data_in[108]
  PIN data_in[109]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.126000 ;
    ANTENNADIFFAREA 0.434700 ;
    PORT
      LAYER met3 ;
        RECT 575.150 365.880 579.150 366.480 ;
    END
  END data_in[109]
  PIN data_in[10]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.126000 ;
    ANTENNADIFFAREA 0.434700 ;
    PORT
      LAYER met3 ;
        RECT 575.150 96.600 579.150 97.200 ;
    END
  END data_in[10]
  PIN data_in[110]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.126000 ;
    ANTENNADIFFAREA 0.434700 ;
    PORT
      LAYER met3 ;
        RECT 575.150 368.600 579.150 369.200 ;
    END
  END data_in[110]
  PIN data_in[111]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.126000 ;
    ANTENNADIFFAREA 0.434700 ;
    PORT
      LAYER met3 ;
        RECT 575.150 371.320 579.150 371.920 ;
    END
  END data_in[111]
  PIN data_in[112]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.126000 ;
    ANTENNADIFFAREA 0.434700 ;
    PORT
      LAYER met3 ;
        RECT 575.150 374.040 579.150 374.640 ;
    END
  END data_in[112]
  PIN data_in[113]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.126000 ;
    ANTENNADIFFAREA 0.434700 ;
    PORT
      LAYER met3 ;
        RECT 575.150 376.760 579.150 377.360 ;
    END
  END data_in[113]
  PIN data_in[114]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.126000 ;
    ANTENNADIFFAREA 0.434700 ;
    PORT
      LAYER met3 ;
        RECT 575.150 379.480 579.150 380.080 ;
    END
  END data_in[114]
  PIN data_in[115]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.126000 ;
    ANTENNADIFFAREA 0.434700 ;
    PORT
      LAYER met3 ;
        RECT 575.150 382.200 579.150 382.800 ;
    END
  END data_in[115]
  PIN data_in[116]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.126000 ;
    ANTENNADIFFAREA 0.434700 ;
    PORT
      LAYER met3 ;
        RECT 575.150 384.920 579.150 385.520 ;
    END
  END data_in[116]
  PIN data_in[117]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.126000 ;
    ANTENNADIFFAREA 0.434700 ;
    PORT
      LAYER met3 ;
        RECT 575.150 387.640 579.150 388.240 ;
    END
  END data_in[117]
  PIN data_in[118]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.126000 ;
    ANTENNADIFFAREA 0.434700 ;
    PORT
      LAYER met3 ;
        RECT 575.150 390.360 579.150 390.960 ;
    END
  END data_in[118]
  PIN data_in[119]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.126000 ;
    ANTENNADIFFAREA 0.434700 ;
    PORT
      LAYER met3 ;
        RECT 575.150 393.080 579.150 393.680 ;
    END
  END data_in[119]
  PIN data_in[11]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.126000 ;
    ANTENNADIFFAREA 0.434700 ;
    PORT
      LAYER met3 ;
        RECT 575.150 99.320 579.150 99.920 ;
    END
  END data_in[11]
  PIN data_in[120]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.126000 ;
    ANTENNADIFFAREA 0.434700 ;
    PORT
      LAYER met3 ;
        RECT 575.150 395.800 579.150 396.400 ;
    END
  END data_in[120]
  PIN data_in[121]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.126000 ;
    ANTENNADIFFAREA 0.434700 ;
    PORT
      LAYER met3 ;
        RECT 575.150 398.520 579.150 399.120 ;
    END
  END data_in[121]
  PIN data_in[122]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.126000 ;
    ANTENNADIFFAREA 0.434700 ;
    PORT
      LAYER met3 ;
        RECT 575.150 401.240 579.150 401.840 ;
    END
  END data_in[122]
  PIN data_in[123]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.126000 ;
    ANTENNADIFFAREA 0.434700 ;
    PORT
      LAYER met3 ;
        RECT 575.150 403.960 579.150 404.560 ;
    END
  END data_in[123]
  PIN data_in[124]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.126000 ;
    ANTENNADIFFAREA 0.434700 ;
    PORT
      LAYER met3 ;
        RECT 575.150 406.680 579.150 407.280 ;
    END
  END data_in[124]
  PIN data_in[125]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.126000 ;
    ANTENNADIFFAREA 0.434700 ;
    PORT
      LAYER met3 ;
        RECT 575.150 409.400 579.150 410.000 ;
    END
  END data_in[125]
  PIN data_in[126]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.126000 ;
    ANTENNADIFFAREA 0.434700 ;
    PORT
      LAYER met3 ;
        RECT 575.150 412.120 579.150 412.720 ;
    END
  END data_in[126]
  PIN data_in[127]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.126000 ;
    ANTENNADIFFAREA 0.434700 ;
    PORT
      LAYER met3 ;
        RECT 575.150 414.840 579.150 415.440 ;
    END
  END data_in[127]
  PIN data_in[128]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.126000 ;
    ANTENNADIFFAREA 0.434700 ;
    PORT
      LAYER met3 ;
        RECT 575.150 417.560 579.150 418.160 ;
    END
  END data_in[128]
  PIN data_in[129]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.126000 ;
    ANTENNADIFFAREA 0.434700 ;
    PORT
      LAYER met3 ;
        RECT 575.150 420.280 579.150 420.880 ;
    END
  END data_in[129]
  PIN data_in[12]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.126000 ;
    ANTENNADIFFAREA 0.434700 ;
    PORT
      LAYER met3 ;
        RECT 575.150 102.040 579.150 102.640 ;
    END
  END data_in[12]
  PIN data_in[130]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.126000 ;
    ANTENNADIFFAREA 0.434700 ;
    PORT
      LAYER met3 ;
        RECT 575.150 423.000 579.150 423.600 ;
    END
  END data_in[130]
  PIN data_in[131]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.126000 ;
    ANTENNADIFFAREA 0.434700 ;
    PORT
      LAYER met3 ;
        RECT 575.150 425.720 579.150 426.320 ;
    END
  END data_in[131]
  PIN data_in[132]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.126000 ;
    ANTENNADIFFAREA 0.434700 ;
    PORT
      LAYER met3 ;
        RECT 575.150 428.440 579.150 429.040 ;
    END
  END data_in[132]
  PIN data_in[133]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.126000 ;
    ANTENNADIFFAREA 0.434700 ;
    PORT
      LAYER met3 ;
        RECT 575.150 431.160 579.150 431.760 ;
    END
  END data_in[133]
  PIN data_in[134]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.126000 ;
    ANTENNADIFFAREA 0.434700 ;
    PORT
      LAYER met3 ;
        RECT 575.150 433.880 579.150 434.480 ;
    END
  END data_in[134]
  PIN data_in[135]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.126000 ;
    ANTENNADIFFAREA 0.434700 ;
    PORT
      LAYER met3 ;
        RECT 575.150 436.600 579.150 437.200 ;
    END
  END data_in[135]
  PIN data_in[136]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.126000 ;
    ANTENNADIFFAREA 0.434700 ;
    PORT
      LAYER met3 ;
        RECT 575.150 439.320 579.150 439.920 ;
    END
  END data_in[136]
  PIN data_in[137]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.126000 ;
    ANTENNADIFFAREA 0.434700 ;
    PORT
      LAYER met3 ;
        RECT 575.150 442.040 579.150 442.640 ;
    END
  END data_in[137]
  PIN data_in[138]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.126000 ;
    ANTENNADIFFAREA 0.434700 ;
    PORT
      LAYER met3 ;
        RECT 575.150 444.760 579.150 445.360 ;
    END
  END data_in[138]
  PIN data_in[139]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.126000 ;
    ANTENNADIFFAREA 0.434700 ;
    PORT
      LAYER met3 ;
        RECT 575.150 447.480 579.150 448.080 ;
    END
  END data_in[139]
  PIN data_in[13]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.126000 ;
    ANTENNADIFFAREA 0.434700 ;
    PORT
      LAYER met3 ;
        RECT 575.150 104.760 579.150 105.360 ;
    END
  END data_in[13]
  PIN data_in[140]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.126000 ;
    ANTENNADIFFAREA 0.434700 ;
    PORT
      LAYER met3 ;
        RECT 575.150 450.200 579.150 450.800 ;
    END
  END data_in[140]
  PIN data_in[141]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.126000 ;
    ANTENNADIFFAREA 0.434700 ;
    PORT
      LAYER met3 ;
        RECT 575.150 452.920 579.150 453.520 ;
    END
  END data_in[141]
  PIN data_in[142]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.126000 ;
    ANTENNADIFFAREA 0.434700 ;
    PORT
      LAYER met3 ;
        RECT 575.150 455.640 579.150 456.240 ;
    END
  END data_in[142]
  PIN data_in[143]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.126000 ;
    ANTENNADIFFAREA 0.434700 ;
    PORT
      LAYER met3 ;
        RECT 575.150 458.360 579.150 458.960 ;
    END
  END data_in[143]
  PIN data_in[144]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.126000 ;
    ANTENNADIFFAREA 0.434700 ;
    PORT
      LAYER met3 ;
        RECT 575.150 461.080 579.150 461.680 ;
    END
  END data_in[144]
  PIN data_in[145]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.126000 ;
    ANTENNADIFFAREA 0.434700 ;
    PORT
      LAYER met3 ;
        RECT 575.150 463.800 579.150 464.400 ;
    END
  END data_in[145]
  PIN data_in[146]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.126000 ;
    ANTENNADIFFAREA 0.434700 ;
    PORT
      LAYER met3 ;
        RECT 575.150 466.520 579.150 467.120 ;
    END
  END data_in[146]
  PIN data_in[147]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.126000 ;
    ANTENNADIFFAREA 0.434700 ;
    PORT
      LAYER met3 ;
        RECT 575.150 469.240 579.150 469.840 ;
    END
  END data_in[147]
  PIN data_in[148]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.126000 ;
    ANTENNADIFFAREA 0.434700 ;
    PORT
      LAYER met3 ;
        RECT 575.150 471.960 579.150 472.560 ;
    END
  END data_in[148]
  PIN data_in[149]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.126000 ;
    ANTENNADIFFAREA 0.434700 ;
    PORT
      LAYER met3 ;
        RECT 575.150 474.680 579.150 475.280 ;
    END
  END data_in[149]
  PIN data_in[14]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.126000 ;
    ANTENNADIFFAREA 0.434700 ;
    PORT
      LAYER met3 ;
        RECT 575.150 107.480 579.150 108.080 ;
    END
  END data_in[14]
  PIN data_in[150]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.126000 ;
    ANTENNADIFFAREA 0.434700 ;
    PORT
      LAYER met3 ;
        RECT 575.150 477.400 579.150 478.000 ;
    END
  END data_in[150]
  PIN data_in[151]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.126000 ;
    ANTENNADIFFAREA 0.434700 ;
    PORT
      LAYER met3 ;
        RECT 575.150 480.120 579.150 480.720 ;
    END
  END data_in[151]
  PIN data_in[152]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.126000 ;
    ANTENNADIFFAREA 0.434700 ;
    PORT
      LAYER met3 ;
        RECT 575.150 482.840 579.150 483.440 ;
    END
  END data_in[152]
  PIN data_in[153]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.126000 ;
    ANTENNADIFFAREA 0.434700 ;
    PORT
      LAYER met3 ;
        RECT 575.150 485.560 579.150 486.160 ;
    END
  END data_in[153]
  PIN data_in[154]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.126000 ;
    ANTENNADIFFAREA 0.434700 ;
    PORT
      LAYER met3 ;
        RECT 575.150 488.280 579.150 488.880 ;
    END
  END data_in[154]
  PIN data_in[155]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.126000 ;
    ANTENNADIFFAREA 0.434700 ;
    PORT
      LAYER met3 ;
        RECT 575.150 491.000 579.150 491.600 ;
    END
  END data_in[155]
  PIN data_in[156]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.126000 ;
    ANTENNADIFFAREA 0.434700 ;
    PORT
      LAYER met3 ;
        RECT 575.150 493.720 579.150 494.320 ;
    END
  END data_in[156]
  PIN data_in[157]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.126000 ;
    ANTENNADIFFAREA 0.434700 ;
    PORT
      LAYER met3 ;
        RECT 575.150 496.440 579.150 497.040 ;
    END
  END data_in[157]
  PIN data_in[158]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.126000 ;
    ANTENNADIFFAREA 0.434700 ;
    PORT
      LAYER met3 ;
        RECT 575.150 499.160 579.150 499.760 ;
    END
  END data_in[158]
  PIN data_in[159]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.126000 ;
    ANTENNADIFFAREA 0.434700 ;
    PORT
      LAYER met3 ;
        RECT 575.150 501.880 579.150 502.480 ;
    END
  END data_in[159]
  PIN data_in[15]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.126000 ;
    ANTENNADIFFAREA 0.434700 ;
    PORT
      LAYER met3 ;
        RECT 575.150 110.200 579.150 110.800 ;
    END
  END data_in[15]
  PIN data_in[160]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.126000 ;
    ANTENNADIFFAREA 0.434700 ;
    PORT
      LAYER met3 ;
        RECT 575.150 504.600 579.150 505.200 ;
    END
  END data_in[160]
  PIN data_in[161]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.126000 ;
    ANTENNADIFFAREA 0.434700 ;
    PORT
      LAYER met3 ;
        RECT 575.150 507.320 579.150 507.920 ;
    END
  END data_in[161]
  PIN data_in[162]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.126000 ;
    ANTENNADIFFAREA 0.434700 ;
    PORT
      LAYER met3 ;
        RECT 575.150 510.040 579.150 510.640 ;
    END
  END data_in[162]
  PIN data_in[16]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.126000 ;
    ANTENNADIFFAREA 0.434700 ;
    PORT
      LAYER met3 ;
        RECT 575.150 112.920 579.150 113.520 ;
    END
  END data_in[16]
  PIN data_in[17]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.126000 ;
    ANTENNADIFFAREA 0.434700 ;
    PORT
      LAYER met3 ;
        RECT 575.150 115.640 579.150 116.240 ;
    END
  END data_in[17]
  PIN data_in[18]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.126000 ;
    ANTENNADIFFAREA 0.434700 ;
    PORT
      LAYER met3 ;
        RECT 575.150 118.360 579.150 118.960 ;
    END
  END data_in[18]
  PIN data_in[19]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.126000 ;
    ANTENNADIFFAREA 0.434700 ;
    PORT
      LAYER met3 ;
        RECT 575.150 121.080 579.150 121.680 ;
    END
  END data_in[19]
  PIN data_in[1]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.126000 ;
    ANTENNADIFFAREA 0.434700 ;
    PORT
      LAYER met3 ;
        RECT 575.150 72.120 579.150 72.720 ;
    END
  END data_in[1]
  PIN data_in[20]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.126000 ;
    ANTENNADIFFAREA 0.434700 ;
    PORT
      LAYER met3 ;
        RECT 575.150 123.800 579.150 124.400 ;
    END
  END data_in[20]
  PIN data_in[21]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.126000 ;
    ANTENNADIFFAREA 0.434700 ;
    PORT
      LAYER met3 ;
        RECT 575.150 126.520 579.150 127.120 ;
    END
  END data_in[21]
  PIN data_in[22]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.126000 ;
    ANTENNADIFFAREA 0.434700 ;
    PORT
      LAYER met3 ;
        RECT 575.150 129.240 579.150 129.840 ;
    END
  END data_in[22]
  PIN data_in[23]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.126000 ;
    ANTENNADIFFAREA 0.434700 ;
    PORT
      LAYER met3 ;
        RECT 575.150 131.960 579.150 132.560 ;
    END
  END data_in[23]
  PIN data_in[24]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.126000 ;
    ANTENNADIFFAREA 0.434700 ;
    PORT
      LAYER met3 ;
        RECT 575.150 134.680 579.150 135.280 ;
    END
  END data_in[24]
  PIN data_in[25]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.126000 ;
    ANTENNADIFFAREA 0.434700 ;
    PORT
      LAYER met3 ;
        RECT 575.150 137.400 579.150 138.000 ;
    END
  END data_in[25]
  PIN data_in[26]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.126000 ;
    ANTENNADIFFAREA 0.434700 ;
    PORT
      LAYER met3 ;
        RECT 575.150 140.120 579.150 140.720 ;
    END
  END data_in[26]
  PIN data_in[27]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.126000 ;
    ANTENNADIFFAREA 0.434700 ;
    PORT
      LAYER met3 ;
        RECT 575.150 142.840 579.150 143.440 ;
    END
  END data_in[27]
  PIN data_in[28]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.126000 ;
    ANTENNADIFFAREA 0.434700 ;
    PORT
      LAYER met3 ;
        RECT 575.150 145.560 579.150 146.160 ;
    END
  END data_in[28]
  PIN data_in[29]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.126000 ;
    ANTENNADIFFAREA 0.434700 ;
    PORT
      LAYER met3 ;
        RECT 575.150 148.280 579.150 148.880 ;
    END
  END data_in[29]
  PIN data_in[2]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.126000 ;
    ANTENNADIFFAREA 0.434700 ;
    PORT
      LAYER met3 ;
        RECT 575.150 74.840 579.150 75.440 ;
    END
  END data_in[2]
  PIN data_in[30]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.126000 ;
    ANTENNADIFFAREA 0.434700 ;
    PORT
      LAYER met3 ;
        RECT 575.150 151.000 579.150 151.600 ;
    END
  END data_in[30]
  PIN data_in[31]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.126000 ;
    ANTENNADIFFAREA 0.434700 ;
    PORT
      LAYER met3 ;
        RECT 575.150 153.720 579.150 154.320 ;
    END
  END data_in[31]
  PIN data_in[32]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.126000 ;
    ANTENNADIFFAREA 0.434700 ;
    PORT
      LAYER met3 ;
        RECT 575.150 156.440 579.150 157.040 ;
    END
  END data_in[32]
  PIN data_in[33]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.126000 ;
    ANTENNADIFFAREA 0.869400 ;
    PORT
      LAYER met3 ;
        RECT 575.150 159.160 579.150 159.760 ;
    END
  END data_in[33]
  PIN data_in[34]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.126000 ;
    ANTENNADIFFAREA 0.434700 ;
    PORT
      LAYER met3 ;
        RECT 575.150 161.880 579.150 162.480 ;
    END
  END data_in[34]
  PIN data_in[35]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.126000 ;
    ANTENNADIFFAREA 0.434700 ;
    PORT
      LAYER met3 ;
        RECT 575.150 164.600 579.150 165.200 ;
    END
  END data_in[35]
  PIN data_in[36]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.126000 ;
    ANTENNADIFFAREA 0.434700 ;
    PORT
      LAYER met3 ;
        RECT 575.150 167.320 579.150 167.920 ;
    END
  END data_in[36]
  PIN data_in[37]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.126000 ;
    ANTENNADIFFAREA 0.434700 ;
    PORT
      LAYER met3 ;
        RECT 575.150 170.040 579.150 170.640 ;
    END
  END data_in[37]
  PIN data_in[38]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.126000 ;
    ANTENNADIFFAREA 0.434700 ;
    PORT
      LAYER met3 ;
        RECT 575.150 172.760 579.150 173.360 ;
    END
  END data_in[38]
  PIN data_in[39]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.126000 ;
    ANTENNADIFFAREA 0.434700 ;
    PORT
      LAYER met3 ;
        RECT 575.150 175.480 579.150 176.080 ;
    END
  END data_in[39]
  PIN data_in[3]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.126000 ;
    ANTENNADIFFAREA 0.434700 ;
    PORT
      LAYER met3 ;
        RECT 575.150 77.560 579.150 78.160 ;
    END
  END data_in[3]
  PIN data_in[40]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.126000 ;
    ANTENNADIFFAREA 0.434700 ;
    PORT
      LAYER met3 ;
        RECT 575.150 178.200 579.150 178.800 ;
    END
  END data_in[40]
  PIN data_in[41]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.126000 ;
    ANTENNADIFFAREA 0.434700 ;
    PORT
      LAYER met3 ;
        RECT 575.150 180.920 579.150 181.520 ;
    END
  END data_in[41]
  PIN data_in[42]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.126000 ;
    ANTENNADIFFAREA 0.434700 ;
    PORT
      LAYER met3 ;
        RECT 575.150 183.640 579.150 184.240 ;
    END
  END data_in[42]
  PIN data_in[43]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.126000 ;
    ANTENNADIFFAREA 0.434700 ;
    PORT
      LAYER met3 ;
        RECT 575.150 186.360 579.150 186.960 ;
    END
  END data_in[43]
  PIN data_in[44]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.126000 ;
    ANTENNADIFFAREA 0.434700 ;
    PORT
      LAYER met3 ;
        RECT 575.150 189.080 579.150 189.680 ;
    END
  END data_in[44]
  PIN data_in[45]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.126000 ;
    ANTENNADIFFAREA 0.434700 ;
    PORT
      LAYER met3 ;
        RECT 575.150 191.800 579.150 192.400 ;
    END
  END data_in[45]
  PIN data_in[46]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.126000 ;
    ANTENNADIFFAREA 0.434700 ;
    PORT
      LAYER met3 ;
        RECT 575.150 194.520 579.150 195.120 ;
    END
  END data_in[46]
  PIN data_in[47]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.126000 ;
    ANTENNADIFFAREA 0.434700 ;
    PORT
      LAYER met3 ;
        RECT 575.150 197.240 579.150 197.840 ;
    END
  END data_in[47]
  PIN data_in[48]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.126000 ;
    ANTENNADIFFAREA 0.434700 ;
    PORT
      LAYER met3 ;
        RECT 575.150 199.960 579.150 200.560 ;
    END
  END data_in[48]
  PIN data_in[49]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.126000 ;
    ANTENNADIFFAREA 0.434700 ;
    PORT
      LAYER met3 ;
        RECT 575.150 202.680 579.150 203.280 ;
    END
  END data_in[49]
  PIN data_in[4]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.126000 ;
    ANTENNADIFFAREA 0.434700 ;
    PORT
      LAYER met3 ;
        RECT 575.150 80.280 579.150 80.880 ;
    END
  END data_in[4]
  PIN data_in[50]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.126000 ;
    ANTENNADIFFAREA 0.434700 ;
    PORT
      LAYER met3 ;
        RECT 575.150 205.400 579.150 206.000 ;
    END
  END data_in[50]
  PIN data_in[51]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.126000 ;
    ANTENNADIFFAREA 0.434700 ;
    PORT
      LAYER met3 ;
        RECT 575.150 208.120 579.150 208.720 ;
    END
  END data_in[51]
  PIN data_in[52]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.126000 ;
    ANTENNADIFFAREA 0.434700 ;
    PORT
      LAYER met3 ;
        RECT 575.150 210.840 579.150 211.440 ;
    END
  END data_in[52]
  PIN data_in[53]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.126000 ;
    ANTENNADIFFAREA 0.434700 ;
    PORT
      LAYER met3 ;
        RECT 575.150 213.560 579.150 214.160 ;
    END
  END data_in[53]
  PIN data_in[54]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.126000 ;
    ANTENNADIFFAREA 0.434700 ;
    PORT
      LAYER met3 ;
        RECT 575.150 216.280 579.150 216.880 ;
    END
  END data_in[54]
  PIN data_in[55]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.126000 ;
    ANTENNADIFFAREA 0.434700 ;
    PORT
      LAYER met3 ;
        RECT 575.150 219.000 579.150 219.600 ;
    END
  END data_in[55]
  PIN data_in[56]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.126000 ;
    ANTENNADIFFAREA 0.434700 ;
    PORT
      LAYER met3 ;
        RECT 575.150 221.720 579.150 222.320 ;
    END
  END data_in[56]
  PIN data_in[57]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.126000 ;
    ANTENNADIFFAREA 0.434700 ;
    PORT
      LAYER met3 ;
        RECT 575.150 224.440 579.150 225.040 ;
    END
  END data_in[57]
  PIN data_in[58]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.126000 ;
    ANTENNADIFFAREA 0.434700 ;
    PORT
      LAYER met3 ;
        RECT 575.150 227.160 579.150 227.760 ;
    END
  END data_in[58]
  PIN data_in[59]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.126000 ;
    ANTENNADIFFAREA 0.434700 ;
    PORT
      LAYER met3 ;
        RECT 575.150 229.880 579.150 230.480 ;
    END
  END data_in[59]
  PIN data_in[5]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.126000 ;
    ANTENNADIFFAREA 0.434700 ;
    PORT
      LAYER met3 ;
        RECT 575.150 83.000 579.150 83.600 ;
    END
  END data_in[5]
  PIN data_in[60]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.126000 ;
    ANTENNADIFFAREA 0.434700 ;
    PORT
      LAYER met3 ;
        RECT 575.150 232.600 579.150 233.200 ;
    END
  END data_in[60]
  PIN data_in[61]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.126000 ;
    ANTENNADIFFAREA 0.434700 ;
    PORT
      LAYER met3 ;
        RECT 575.150 235.320 579.150 235.920 ;
    END
  END data_in[61]
  PIN data_in[62]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.126000 ;
    ANTENNADIFFAREA 0.434700 ;
    PORT
      LAYER met3 ;
        RECT 575.150 238.040 579.150 238.640 ;
    END
  END data_in[62]
  PIN data_in[63]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.126000 ;
    ANTENNADIFFAREA 0.434700 ;
    PORT
      LAYER met3 ;
        RECT 575.150 240.760 579.150 241.360 ;
    END
  END data_in[63]
  PIN data_in[64]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.126000 ;
    ANTENNADIFFAREA 0.434700 ;
    PORT
      LAYER met3 ;
        RECT 575.150 243.480 579.150 244.080 ;
    END
  END data_in[64]
  PIN data_in[65]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.126000 ;
    ANTENNADIFFAREA 0.434700 ;
    PORT
      LAYER met3 ;
        RECT 575.150 246.200 579.150 246.800 ;
    END
  END data_in[65]
  PIN data_in[66]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.126000 ;
    ANTENNADIFFAREA 0.434700 ;
    PORT
      LAYER met3 ;
        RECT 575.150 248.920 579.150 249.520 ;
    END
  END data_in[66]
  PIN data_in[67]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.126000 ;
    ANTENNADIFFAREA 0.434700 ;
    PORT
      LAYER met3 ;
        RECT 575.150 251.640 579.150 252.240 ;
    END
  END data_in[67]
  PIN data_in[68]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.126000 ;
    ANTENNADIFFAREA 0.434700 ;
    PORT
      LAYER met3 ;
        RECT 575.150 254.360 579.150 254.960 ;
    END
  END data_in[68]
  PIN data_in[69]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.126000 ;
    ANTENNADIFFAREA 0.434700 ;
    PORT
      LAYER met3 ;
        RECT 575.150 257.080 579.150 257.680 ;
    END
  END data_in[69]
  PIN data_in[6]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.126000 ;
    ANTENNADIFFAREA 0.434700 ;
    PORT
      LAYER met3 ;
        RECT 575.150 85.720 579.150 86.320 ;
    END
  END data_in[6]
  PIN data_in[70]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.126000 ;
    ANTENNADIFFAREA 0.434700 ;
    PORT
      LAYER met3 ;
        RECT 575.150 259.800 579.150 260.400 ;
    END
  END data_in[70]
  PIN data_in[71]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.126000 ;
    ANTENNADIFFAREA 0.434700 ;
    PORT
      LAYER met3 ;
        RECT 575.150 262.520 579.150 263.120 ;
    END
  END data_in[71]
  PIN data_in[72]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.126000 ;
    ANTENNADIFFAREA 0.434700 ;
    PORT
      LAYER met3 ;
        RECT 575.150 265.240 579.150 265.840 ;
    END
  END data_in[72]
  PIN data_in[73]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.126000 ;
    ANTENNADIFFAREA 0.434700 ;
    PORT
      LAYER met3 ;
        RECT 575.150 267.960 579.150 268.560 ;
    END
  END data_in[73]
  PIN data_in[74]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.126000 ;
    ANTENNADIFFAREA 0.434700 ;
    PORT
      LAYER met3 ;
        RECT 575.150 270.680 579.150 271.280 ;
    END
  END data_in[74]
  PIN data_in[75]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.126000 ;
    ANTENNADIFFAREA 0.434700 ;
    PORT
      LAYER met3 ;
        RECT 575.150 273.400 579.150 274.000 ;
    END
  END data_in[75]
  PIN data_in[76]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.126000 ;
    ANTENNADIFFAREA 0.434700 ;
    PORT
      LAYER met3 ;
        RECT 575.150 276.120 579.150 276.720 ;
    END
  END data_in[76]
  PIN data_in[77]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.126000 ;
    ANTENNADIFFAREA 0.434700 ;
    PORT
      LAYER met3 ;
        RECT 575.150 278.840 579.150 279.440 ;
    END
  END data_in[77]
  PIN data_in[78]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.126000 ;
    ANTENNADIFFAREA 0.434700 ;
    PORT
      LAYER met3 ;
        RECT 575.150 281.560 579.150 282.160 ;
    END
  END data_in[78]
  PIN data_in[79]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.126000 ;
    ANTENNADIFFAREA 0.434700 ;
    PORT
      LAYER met3 ;
        RECT 575.150 284.280 579.150 284.880 ;
    END
  END data_in[79]
  PIN data_in[7]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.126000 ;
    ANTENNADIFFAREA 0.434700 ;
    PORT
      LAYER met3 ;
        RECT 575.150 88.440 579.150 89.040 ;
    END
  END data_in[7]
  PIN data_in[80]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.126000 ;
    ANTENNADIFFAREA 0.434700 ;
    PORT
      LAYER met3 ;
        RECT 575.150 287.000 579.150 287.600 ;
    END
  END data_in[80]
  PIN data_in[81]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.126000 ;
    ANTENNADIFFAREA 0.434700 ;
    PORT
      LAYER met3 ;
        RECT 575.150 289.720 579.150 290.320 ;
    END
  END data_in[81]
  PIN data_in[82]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.126000 ;
    ANTENNADIFFAREA 0.869400 ;
    PORT
      LAYER met3 ;
        RECT 575.150 292.440 579.150 293.040 ;
    END
  END data_in[82]
  PIN data_in[83]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.126000 ;
    ANTENNADIFFAREA 0.434700 ;
    PORT
      LAYER met3 ;
        RECT 575.150 295.160 579.150 295.760 ;
    END
  END data_in[83]
  PIN data_in[84]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.126000 ;
    ANTENNADIFFAREA 0.434700 ;
    PORT
      LAYER met3 ;
        RECT 575.150 297.880 579.150 298.480 ;
    END
  END data_in[84]
  PIN data_in[85]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.126000 ;
    ANTENNADIFFAREA 0.434700 ;
    PORT
      LAYER met3 ;
        RECT 575.150 300.600 579.150 301.200 ;
    END
  END data_in[85]
  PIN data_in[86]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.126000 ;
    ANTENNADIFFAREA 0.434700 ;
    PORT
      LAYER met3 ;
        RECT 575.150 303.320 579.150 303.920 ;
    END
  END data_in[86]
  PIN data_in[87]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.126000 ;
    ANTENNADIFFAREA 0.434700 ;
    PORT
      LAYER met3 ;
        RECT 575.150 306.040 579.150 306.640 ;
    END
  END data_in[87]
  PIN data_in[88]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.126000 ;
    ANTENNADIFFAREA 0.434700 ;
    PORT
      LAYER met3 ;
        RECT 575.150 308.760 579.150 309.360 ;
    END
  END data_in[88]
  PIN data_in[89]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.126000 ;
    ANTENNADIFFAREA 0.434700 ;
    PORT
      LAYER met3 ;
        RECT 575.150 311.480 579.150 312.080 ;
    END
  END data_in[89]
  PIN data_in[8]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.126000 ;
    ANTENNADIFFAREA 0.434700 ;
    PORT
      LAYER met3 ;
        RECT 575.150 91.160 579.150 91.760 ;
    END
  END data_in[8]
  PIN data_in[90]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.126000 ;
    ANTENNADIFFAREA 0.434700 ;
    PORT
      LAYER met3 ;
        RECT 575.150 314.200 579.150 314.800 ;
    END
  END data_in[90]
  PIN data_in[91]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.126000 ;
    ANTENNADIFFAREA 0.434700 ;
    PORT
      LAYER met3 ;
        RECT 575.150 316.920 579.150 317.520 ;
    END
  END data_in[91]
  PIN data_in[92]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.126000 ;
    ANTENNADIFFAREA 0.434700 ;
    PORT
      LAYER met3 ;
        RECT 575.150 319.640 579.150 320.240 ;
    END
  END data_in[92]
  PIN data_in[93]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.126000 ;
    ANTENNADIFFAREA 0.434700 ;
    PORT
      LAYER met3 ;
        RECT 575.150 322.360 579.150 322.960 ;
    END
  END data_in[93]
  PIN data_in[94]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.126000 ;
    ANTENNADIFFAREA 0.434700 ;
    PORT
      LAYER met3 ;
        RECT 575.150 325.080 579.150 325.680 ;
    END
  END data_in[94]
  PIN data_in[95]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.126000 ;
    ANTENNADIFFAREA 0.434700 ;
    PORT
      LAYER met3 ;
        RECT 575.150 327.800 579.150 328.400 ;
    END
  END data_in[95]
  PIN data_in[96]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.126000 ;
    ANTENNADIFFAREA 0.434700 ;
    PORT
      LAYER met3 ;
        RECT 575.150 330.520 579.150 331.120 ;
    END
  END data_in[96]
  PIN data_in[97]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.126000 ;
    ANTENNADIFFAREA 0.434700 ;
    PORT
      LAYER met3 ;
        RECT 575.150 333.240 579.150 333.840 ;
    END
  END data_in[97]
  PIN data_in[98]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.126000 ;
    ANTENNADIFFAREA 0.434700 ;
    PORT
      LAYER met3 ;
        RECT 575.150 335.960 579.150 336.560 ;
    END
  END data_in[98]
  PIN data_in[99]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.126000 ;
    ANTENNADIFFAREA 0.434700 ;
    PORT
      LAYER met3 ;
        RECT 575.150 338.680 579.150 339.280 ;
    END
  END data_in[99]
  PIN data_in[9]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.126000 ;
    ANTENNADIFFAREA 0.434700 ;
    PORT
      LAYER met3 ;
        RECT 575.150 93.880 579.150 94.480 ;
    END
  END data_in[9]
  PIN data_out[0]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 2.673000 ;
    PORT
      LAYER met3 ;
        RECT 0.000 68.040 4.000 68.640 ;
    END
  END data_out[0]
  PIN data_out[100]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 2.673000 ;
    PORT
      LAYER met3 ;
        RECT 0.000 340.040 4.000 340.640 ;
    END
  END data_out[100]
  PIN data_out[101]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 2.673000 ;
    PORT
      LAYER met3 ;
        RECT 0.000 342.760 4.000 343.360 ;
    END
  END data_out[101]
  PIN data_out[102]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 2.673000 ;
    PORT
      LAYER met3 ;
        RECT 0.000 345.480 4.000 346.080 ;
    END
  END data_out[102]
  PIN data_out[103]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 2.673000 ;
    PORT
      LAYER met3 ;
        RECT 0.000 348.200 4.000 348.800 ;
    END
  END data_out[103]
  PIN data_out[104]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 2.673000 ;
    PORT
      LAYER met3 ;
        RECT 0.000 350.920 4.000 351.520 ;
    END
  END data_out[104]
  PIN data_out[105]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 2.673000 ;
    PORT
      LAYER met3 ;
        RECT 0.000 353.640 4.000 354.240 ;
    END
  END data_out[105]
  PIN data_out[106]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 2.673000 ;
    PORT
      LAYER met3 ;
        RECT 0.000 356.360 4.000 356.960 ;
    END
  END data_out[106]
  PIN data_out[107]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 2.673000 ;
    PORT
      LAYER met3 ;
        RECT 0.000 359.080 4.000 359.680 ;
    END
  END data_out[107]
  PIN data_out[108]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 2.673000 ;
    PORT
      LAYER met3 ;
        RECT 0.000 361.800 4.000 362.400 ;
    END
  END data_out[108]
  PIN data_out[109]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 2.673000 ;
    PORT
      LAYER met3 ;
        RECT 0.000 364.520 4.000 365.120 ;
    END
  END data_out[109]
  PIN data_out[10]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 2.673000 ;
    PORT
      LAYER met3 ;
        RECT 0.000 95.240 4.000 95.840 ;
    END
  END data_out[10]
  PIN data_out[110]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 2.673000 ;
    PORT
      LAYER met3 ;
        RECT 0.000 367.240 4.000 367.840 ;
    END
  END data_out[110]
  PIN data_out[111]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 2.673000 ;
    PORT
      LAYER met3 ;
        RECT 0.000 369.960 4.000 370.560 ;
    END
  END data_out[111]
  PIN data_out[112]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 2.673000 ;
    PORT
      LAYER met3 ;
        RECT 0.000 372.680 4.000 373.280 ;
    END
  END data_out[112]
  PIN data_out[113]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 2.673000 ;
    PORT
      LAYER met3 ;
        RECT 0.000 375.400 4.000 376.000 ;
    END
  END data_out[113]
  PIN data_out[114]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 2.673000 ;
    PORT
      LAYER met3 ;
        RECT 0.000 378.120 4.000 378.720 ;
    END
  END data_out[114]
  PIN data_out[115]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 2.673000 ;
    PORT
      LAYER met3 ;
        RECT 0.000 380.840 4.000 381.440 ;
    END
  END data_out[115]
  PIN data_out[116]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 2.673000 ;
    PORT
      LAYER met3 ;
        RECT 0.000 383.560 4.000 384.160 ;
    END
  END data_out[116]
  PIN data_out[117]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 2.673000 ;
    PORT
      LAYER met3 ;
        RECT 0.000 386.280 4.000 386.880 ;
    END
  END data_out[117]
  PIN data_out[118]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 2.673000 ;
    PORT
      LAYER met3 ;
        RECT 0.000 389.000 4.000 389.600 ;
    END
  END data_out[118]
  PIN data_out[119]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 2.673000 ;
    PORT
      LAYER met3 ;
        RECT 0.000 391.720 4.000 392.320 ;
    END
  END data_out[119]
  PIN data_out[11]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 2.673000 ;
    PORT
      LAYER met3 ;
        RECT 0.000 97.960 4.000 98.560 ;
    END
  END data_out[11]
  PIN data_out[120]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 2.673000 ;
    PORT
      LAYER met3 ;
        RECT 0.000 394.440 4.000 395.040 ;
    END
  END data_out[120]
  PIN data_out[121]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 2.673000 ;
    PORT
      LAYER met3 ;
        RECT 0.000 397.160 4.000 397.760 ;
    END
  END data_out[121]
  PIN data_out[122]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 2.673000 ;
    PORT
      LAYER met3 ;
        RECT 0.000 399.880 4.000 400.480 ;
    END
  END data_out[122]
  PIN data_out[123]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 2.673000 ;
    PORT
      LAYER met3 ;
        RECT 0.000 402.600 4.000 403.200 ;
    END
  END data_out[123]
  PIN data_out[124]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 2.673000 ;
    PORT
      LAYER met3 ;
        RECT 0.000 405.320 4.000 405.920 ;
    END
  END data_out[124]
  PIN data_out[125]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 2.673000 ;
    PORT
      LAYER met3 ;
        RECT 0.000 408.040 4.000 408.640 ;
    END
  END data_out[125]
  PIN data_out[126]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 2.673000 ;
    PORT
      LAYER met3 ;
        RECT 0.000 410.760 4.000 411.360 ;
    END
  END data_out[126]
  PIN data_out[127]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 2.673000 ;
    PORT
      LAYER met3 ;
        RECT 0.000 413.480 4.000 414.080 ;
    END
  END data_out[127]
  PIN data_out[128]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 2.673000 ;
    PORT
      LAYER met3 ;
        RECT 0.000 416.200 4.000 416.800 ;
    END
  END data_out[128]
  PIN data_out[129]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 2.673000 ;
    PORT
      LAYER met3 ;
        RECT 0.000 418.920 4.000 419.520 ;
    END
  END data_out[129]
  PIN data_out[12]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 2.673000 ;
    PORT
      LAYER met3 ;
        RECT 0.000 100.680 4.000 101.280 ;
    END
  END data_out[12]
  PIN data_out[130]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 2.673000 ;
    PORT
      LAYER met3 ;
        RECT 0.000 421.640 4.000 422.240 ;
    END
  END data_out[130]
  PIN data_out[131]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 2.673000 ;
    PORT
      LAYER met3 ;
        RECT 0.000 424.360 4.000 424.960 ;
    END
  END data_out[131]
  PIN data_out[132]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 2.673000 ;
    PORT
      LAYER met3 ;
        RECT 0.000 427.080 4.000 427.680 ;
    END
  END data_out[132]
  PIN data_out[133]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 2.673000 ;
    PORT
      LAYER met3 ;
        RECT 0.000 429.800 4.000 430.400 ;
    END
  END data_out[133]
  PIN data_out[134]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 2.673000 ;
    PORT
      LAYER met3 ;
        RECT 0.000 432.520 4.000 433.120 ;
    END
  END data_out[134]
  PIN data_out[135]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 2.673000 ;
    PORT
      LAYER met3 ;
        RECT 0.000 435.240 4.000 435.840 ;
    END
  END data_out[135]
  PIN data_out[136]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 2.673000 ;
    PORT
      LAYER met3 ;
        RECT 0.000 437.960 4.000 438.560 ;
    END
  END data_out[136]
  PIN data_out[137]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 2.673000 ;
    PORT
      LAYER met3 ;
        RECT 0.000 440.680 4.000 441.280 ;
    END
  END data_out[137]
  PIN data_out[138]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 2.673000 ;
    PORT
      LAYER met3 ;
        RECT 0.000 443.400 4.000 444.000 ;
    END
  END data_out[138]
  PIN data_out[139]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 2.673000 ;
    PORT
      LAYER met3 ;
        RECT 0.000 446.120 4.000 446.720 ;
    END
  END data_out[139]
  PIN data_out[13]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 2.673000 ;
    PORT
      LAYER met3 ;
        RECT 0.000 103.400 4.000 104.000 ;
    END
  END data_out[13]
  PIN data_out[140]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 2.673000 ;
    PORT
      LAYER met3 ;
        RECT 0.000 448.840 4.000 449.440 ;
    END
  END data_out[140]
  PIN data_out[141]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 2.673000 ;
    PORT
      LAYER met3 ;
        RECT 0.000 451.560 4.000 452.160 ;
    END
  END data_out[141]
  PIN data_out[142]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 2.673000 ;
    PORT
      LAYER met3 ;
        RECT 0.000 454.280 4.000 454.880 ;
    END
  END data_out[142]
  PIN data_out[143]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 2.673000 ;
    PORT
      LAYER met3 ;
        RECT 0.000 457.000 4.000 457.600 ;
    END
  END data_out[143]
  PIN data_out[144]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 2.673000 ;
    PORT
      LAYER met3 ;
        RECT 0.000 459.720 4.000 460.320 ;
    END
  END data_out[144]
  PIN data_out[145]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 2.673000 ;
    PORT
      LAYER met3 ;
        RECT 0.000 462.440 4.000 463.040 ;
    END
  END data_out[145]
  PIN data_out[146]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 2.673000 ;
    PORT
      LAYER met3 ;
        RECT 0.000 465.160 4.000 465.760 ;
    END
  END data_out[146]
  PIN data_out[147]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 2.673000 ;
    PORT
      LAYER met3 ;
        RECT 0.000 467.880 4.000 468.480 ;
    END
  END data_out[147]
  PIN data_out[148]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 2.673000 ;
    PORT
      LAYER met3 ;
        RECT 0.000 470.600 4.000 471.200 ;
    END
  END data_out[148]
  PIN data_out[149]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 2.673000 ;
    PORT
      LAYER met3 ;
        RECT 0.000 473.320 4.000 473.920 ;
    END
  END data_out[149]
  PIN data_out[14]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 2.673000 ;
    PORT
      LAYER met3 ;
        RECT 0.000 106.120 4.000 106.720 ;
    END
  END data_out[14]
  PIN data_out[150]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 2.673000 ;
    PORT
      LAYER met3 ;
        RECT 0.000 476.040 4.000 476.640 ;
    END
  END data_out[150]
  PIN data_out[151]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 2.673000 ;
    PORT
      LAYER met3 ;
        RECT 0.000 478.760 4.000 479.360 ;
    END
  END data_out[151]
  PIN data_out[152]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 2.673000 ;
    PORT
      LAYER met3 ;
        RECT 0.000 481.480 4.000 482.080 ;
    END
  END data_out[152]
  PIN data_out[153]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 2.673000 ;
    PORT
      LAYER met3 ;
        RECT 0.000 484.200 4.000 484.800 ;
    END
  END data_out[153]
  PIN data_out[154]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 2.673000 ;
    PORT
      LAYER met3 ;
        RECT 0.000 486.920 4.000 487.520 ;
    END
  END data_out[154]
  PIN data_out[155]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 2.673000 ;
    PORT
      LAYER met3 ;
        RECT 0.000 489.640 4.000 490.240 ;
    END
  END data_out[155]
  PIN data_out[156]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 2.673000 ;
    PORT
      LAYER met3 ;
        RECT 0.000 492.360 4.000 492.960 ;
    END
  END data_out[156]
  PIN data_out[157]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 2.673000 ;
    PORT
      LAYER met3 ;
        RECT 0.000 495.080 4.000 495.680 ;
    END
  END data_out[157]
  PIN data_out[158]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 2.673000 ;
    PORT
      LAYER met3 ;
        RECT 0.000 497.800 4.000 498.400 ;
    END
  END data_out[158]
  PIN data_out[159]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 2.673000 ;
    PORT
      LAYER met3 ;
        RECT 0.000 500.520 4.000 501.120 ;
    END
  END data_out[159]
  PIN data_out[15]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 2.673000 ;
    PORT
      LAYER met3 ;
        RECT 0.000 108.840 4.000 109.440 ;
    END
  END data_out[15]
  PIN data_out[160]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 2.673000 ;
    PORT
      LAYER met3 ;
        RECT 0.000 503.240 4.000 503.840 ;
    END
  END data_out[160]
  PIN data_out[161]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 2.673000 ;
    PORT
      LAYER met3 ;
        RECT 0.000 505.960 4.000 506.560 ;
    END
  END data_out[161]
  PIN data_out[162]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 2.673000 ;
    PORT
      LAYER met3 ;
        RECT 0.000 508.680 4.000 509.280 ;
    END
  END data_out[162]
  PIN data_out[16]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 2.673000 ;
    PORT
      LAYER met3 ;
        RECT 0.000 111.560 4.000 112.160 ;
    END
  END data_out[16]
  PIN data_out[17]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 2.673000 ;
    PORT
      LAYER met3 ;
        RECT 0.000 114.280 4.000 114.880 ;
    END
  END data_out[17]
  PIN data_out[18]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 2.673000 ;
    PORT
      LAYER met3 ;
        RECT 0.000 117.000 4.000 117.600 ;
    END
  END data_out[18]
  PIN data_out[19]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 2.673000 ;
    PORT
      LAYER met3 ;
        RECT 0.000 119.720 4.000 120.320 ;
    END
  END data_out[19]
  PIN data_out[1]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 2.673000 ;
    PORT
      LAYER met3 ;
        RECT 0.000 70.760 4.000 71.360 ;
    END
  END data_out[1]
  PIN data_out[20]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 2.673000 ;
    PORT
      LAYER met3 ;
        RECT 0.000 122.440 4.000 123.040 ;
    END
  END data_out[20]
  PIN data_out[21]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 2.673000 ;
    PORT
      LAYER met3 ;
        RECT 0.000 125.160 4.000 125.760 ;
    END
  END data_out[21]
  PIN data_out[22]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 2.673000 ;
    PORT
      LAYER met3 ;
        RECT 0.000 127.880 4.000 128.480 ;
    END
  END data_out[22]
  PIN data_out[23]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 2.673000 ;
    PORT
      LAYER met3 ;
        RECT 0.000 130.600 4.000 131.200 ;
    END
  END data_out[23]
  PIN data_out[24]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 2.673000 ;
    PORT
      LAYER met3 ;
        RECT 0.000 133.320 4.000 133.920 ;
    END
  END data_out[24]
  PIN data_out[25]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 2.673000 ;
    PORT
      LAYER met3 ;
        RECT 0.000 136.040 4.000 136.640 ;
    END
  END data_out[25]
  PIN data_out[26]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 2.673000 ;
    PORT
      LAYER met3 ;
        RECT 0.000 138.760 4.000 139.360 ;
    END
  END data_out[26]
  PIN data_out[27]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 2.673000 ;
    PORT
      LAYER met3 ;
        RECT 0.000 141.480 4.000 142.080 ;
    END
  END data_out[27]
  PIN data_out[28]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 2.673000 ;
    PORT
      LAYER met3 ;
        RECT 0.000 144.200 4.000 144.800 ;
    END
  END data_out[28]
  PIN data_out[29]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 2.673000 ;
    PORT
      LAYER met3 ;
        RECT 0.000 146.920 4.000 147.520 ;
    END
  END data_out[29]
  PIN data_out[2]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 2.673000 ;
    PORT
      LAYER met3 ;
        RECT 0.000 73.480 4.000 74.080 ;
    END
  END data_out[2]
  PIN data_out[30]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 2.673000 ;
    PORT
      LAYER met3 ;
        RECT 0.000 149.640 4.000 150.240 ;
    END
  END data_out[30]
  PIN data_out[31]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 2.673000 ;
    PORT
      LAYER met3 ;
        RECT 0.000 152.360 4.000 152.960 ;
    END
  END data_out[31]
  PIN data_out[32]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 2.673000 ;
    PORT
      LAYER met3 ;
        RECT 0.000 155.080 4.000 155.680 ;
    END
  END data_out[32]
  PIN data_out[33]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 2.673000 ;
    PORT
      LAYER met3 ;
        RECT 0.000 157.800 4.000 158.400 ;
    END
  END data_out[33]
  PIN data_out[34]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 2.673000 ;
    PORT
      LAYER met3 ;
        RECT 0.000 160.520 4.000 161.120 ;
    END
  END data_out[34]
  PIN data_out[35]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 2.673000 ;
    PORT
      LAYER met3 ;
        RECT 0.000 163.240 4.000 163.840 ;
    END
  END data_out[35]
  PIN data_out[36]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 2.673000 ;
    PORT
      LAYER met3 ;
        RECT 0.000 165.960 4.000 166.560 ;
    END
  END data_out[36]
  PIN data_out[37]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 2.673000 ;
    PORT
      LAYER met3 ;
        RECT 0.000 168.680 4.000 169.280 ;
    END
  END data_out[37]
  PIN data_out[38]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 2.673000 ;
    PORT
      LAYER met3 ;
        RECT 0.000 171.400 4.000 172.000 ;
    END
  END data_out[38]
  PIN data_out[39]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 2.673000 ;
    PORT
      LAYER met3 ;
        RECT 0.000 174.120 4.000 174.720 ;
    END
  END data_out[39]
  PIN data_out[3]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 2.673000 ;
    PORT
      LAYER met3 ;
        RECT 0.000 76.200 4.000 76.800 ;
    END
  END data_out[3]
  PIN data_out[40]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 2.673000 ;
    PORT
      LAYER met3 ;
        RECT 0.000 176.840 4.000 177.440 ;
    END
  END data_out[40]
  PIN data_out[41]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 2.673000 ;
    PORT
      LAYER met3 ;
        RECT 0.000 179.560 4.000 180.160 ;
    END
  END data_out[41]
  PIN data_out[42]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 2.673000 ;
    PORT
      LAYER met3 ;
        RECT 0.000 182.280 4.000 182.880 ;
    END
  END data_out[42]
  PIN data_out[43]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 2.673000 ;
    PORT
      LAYER met3 ;
        RECT 0.000 185.000 4.000 185.600 ;
    END
  END data_out[43]
  PIN data_out[44]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 2.673000 ;
    PORT
      LAYER met3 ;
        RECT 0.000 187.720 4.000 188.320 ;
    END
  END data_out[44]
  PIN data_out[45]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 2.673000 ;
    PORT
      LAYER met3 ;
        RECT 0.000 190.440 4.000 191.040 ;
    END
  END data_out[45]
  PIN data_out[46]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 2.673000 ;
    PORT
      LAYER met3 ;
        RECT 0.000 193.160 4.000 193.760 ;
    END
  END data_out[46]
  PIN data_out[47]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 2.673000 ;
    PORT
      LAYER met3 ;
        RECT 0.000 195.880 4.000 196.480 ;
    END
  END data_out[47]
  PIN data_out[48]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 2.673000 ;
    PORT
      LAYER met3 ;
        RECT 0.000 198.600 4.000 199.200 ;
    END
  END data_out[48]
  PIN data_out[49]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 2.673000 ;
    PORT
      LAYER met3 ;
        RECT 0.000 201.320 4.000 201.920 ;
    END
  END data_out[49]
  PIN data_out[4]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 2.673000 ;
    PORT
      LAYER met3 ;
        RECT 0.000 78.920 4.000 79.520 ;
    END
  END data_out[4]
  PIN data_out[50]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 2.673000 ;
    PORT
      LAYER met3 ;
        RECT 0.000 204.040 4.000 204.640 ;
    END
  END data_out[50]
  PIN data_out[51]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 2.673000 ;
    PORT
      LAYER met3 ;
        RECT 0.000 206.760 4.000 207.360 ;
    END
  END data_out[51]
  PIN data_out[52]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 2.673000 ;
    PORT
      LAYER met3 ;
        RECT 0.000 209.480 4.000 210.080 ;
    END
  END data_out[52]
  PIN data_out[53]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 2.673000 ;
    PORT
      LAYER met3 ;
        RECT 0.000 212.200 4.000 212.800 ;
    END
  END data_out[53]
  PIN data_out[54]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 2.673000 ;
    PORT
      LAYER met3 ;
        RECT 0.000 214.920 4.000 215.520 ;
    END
  END data_out[54]
  PIN data_out[55]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 2.673000 ;
    PORT
      LAYER met3 ;
        RECT 0.000 217.640 4.000 218.240 ;
    END
  END data_out[55]
  PIN data_out[56]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 2.673000 ;
    PORT
      LAYER met3 ;
        RECT 0.000 220.360 4.000 220.960 ;
    END
  END data_out[56]
  PIN data_out[57]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 2.673000 ;
    PORT
      LAYER met3 ;
        RECT 0.000 223.080 4.000 223.680 ;
    END
  END data_out[57]
  PIN data_out[58]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 2.673000 ;
    PORT
      LAYER met3 ;
        RECT 0.000 225.800 4.000 226.400 ;
    END
  END data_out[58]
  PIN data_out[59]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 2.673000 ;
    PORT
      LAYER met3 ;
        RECT 0.000 228.520 4.000 229.120 ;
    END
  END data_out[59]
  PIN data_out[5]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 2.673000 ;
    PORT
      LAYER met3 ;
        RECT 0.000 81.640 4.000 82.240 ;
    END
  END data_out[5]
  PIN data_out[60]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 2.673000 ;
    PORT
      LAYER met3 ;
        RECT 0.000 231.240 4.000 231.840 ;
    END
  END data_out[60]
  PIN data_out[61]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 2.673000 ;
    PORT
      LAYER met3 ;
        RECT 0.000 233.960 4.000 234.560 ;
    END
  END data_out[61]
  PIN data_out[62]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 2.673000 ;
    PORT
      LAYER met3 ;
        RECT 0.000 236.680 4.000 237.280 ;
    END
  END data_out[62]
  PIN data_out[63]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 2.673000 ;
    PORT
      LAYER met3 ;
        RECT 0.000 239.400 4.000 240.000 ;
    END
  END data_out[63]
  PIN data_out[64]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 2.673000 ;
    PORT
      LAYER met3 ;
        RECT 0.000 242.120 4.000 242.720 ;
    END
  END data_out[64]
  PIN data_out[65]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 2.673000 ;
    PORT
      LAYER met3 ;
        RECT 0.000 244.840 4.000 245.440 ;
    END
  END data_out[65]
  PIN data_out[66]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 2.673000 ;
    PORT
      LAYER met3 ;
        RECT 0.000 247.560 4.000 248.160 ;
    END
  END data_out[66]
  PIN data_out[67]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 2.673000 ;
    PORT
      LAYER met3 ;
        RECT 0.000 250.280 4.000 250.880 ;
    END
  END data_out[67]
  PIN data_out[68]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 2.673000 ;
    PORT
      LAYER met3 ;
        RECT 0.000 253.000 4.000 253.600 ;
    END
  END data_out[68]
  PIN data_out[69]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 2.673000 ;
    PORT
      LAYER met3 ;
        RECT 0.000 255.720 4.000 256.320 ;
    END
  END data_out[69]
  PIN data_out[6]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 2.673000 ;
    PORT
      LAYER met3 ;
        RECT 0.000 84.360 4.000 84.960 ;
    END
  END data_out[6]
  PIN data_out[70]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 2.673000 ;
    PORT
      LAYER met3 ;
        RECT 0.000 258.440 4.000 259.040 ;
    END
  END data_out[70]
  PIN data_out[71]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 2.673000 ;
    PORT
      LAYER met3 ;
        RECT 0.000 261.160 4.000 261.760 ;
    END
  END data_out[71]
  PIN data_out[72]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 2.673000 ;
    PORT
      LAYER met3 ;
        RECT 0.000 263.880 4.000 264.480 ;
    END
  END data_out[72]
  PIN data_out[73]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 2.673000 ;
    PORT
      LAYER met3 ;
        RECT 0.000 266.600 4.000 267.200 ;
    END
  END data_out[73]
  PIN data_out[74]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 2.673000 ;
    PORT
      LAYER met3 ;
        RECT 0.000 269.320 4.000 269.920 ;
    END
  END data_out[74]
  PIN data_out[75]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 2.673000 ;
    PORT
      LAYER met3 ;
        RECT 0.000 272.040 4.000 272.640 ;
    END
  END data_out[75]
  PIN data_out[76]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 2.673000 ;
    PORT
      LAYER met3 ;
        RECT 0.000 274.760 4.000 275.360 ;
    END
  END data_out[76]
  PIN data_out[77]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 2.673000 ;
    PORT
      LAYER met3 ;
        RECT 0.000 277.480 4.000 278.080 ;
    END
  END data_out[77]
  PIN data_out[78]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 2.673000 ;
    PORT
      LAYER met3 ;
        RECT 0.000 280.200 4.000 280.800 ;
    END
  END data_out[78]
  PIN data_out[79]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 2.673000 ;
    PORT
      LAYER met3 ;
        RECT 0.000 282.920 4.000 283.520 ;
    END
  END data_out[79]
  PIN data_out[7]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 2.673000 ;
    PORT
      LAYER met3 ;
        RECT 0.000 87.080 4.000 87.680 ;
    END
  END data_out[7]
  PIN data_out[80]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 2.673000 ;
    PORT
      LAYER met3 ;
        RECT 0.000 285.640 4.000 286.240 ;
    END
  END data_out[80]
  PIN data_out[81]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 2.673000 ;
    PORT
      LAYER met3 ;
        RECT 0.000 288.360 4.000 288.960 ;
    END
  END data_out[81]
  PIN data_out[82]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 2.673000 ;
    PORT
      LAYER met3 ;
        RECT 0.000 291.080 4.000 291.680 ;
    END
  END data_out[82]
  PIN data_out[83]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 2.673000 ;
    PORT
      LAYER met3 ;
        RECT 0.000 293.800 4.000 294.400 ;
    END
  END data_out[83]
  PIN data_out[84]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 2.673000 ;
    PORT
      LAYER met3 ;
        RECT 0.000 296.520 4.000 297.120 ;
    END
  END data_out[84]
  PIN data_out[85]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 2.673000 ;
    PORT
      LAYER met3 ;
        RECT 0.000 299.240 4.000 299.840 ;
    END
  END data_out[85]
  PIN data_out[86]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 2.673000 ;
    PORT
      LAYER met3 ;
        RECT 0.000 301.960 4.000 302.560 ;
    END
  END data_out[86]
  PIN data_out[87]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 2.673000 ;
    PORT
      LAYER met3 ;
        RECT 0.000 304.680 4.000 305.280 ;
    END
  END data_out[87]
  PIN data_out[88]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 2.673000 ;
    PORT
      LAYER met3 ;
        RECT 0.000 307.400 4.000 308.000 ;
    END
  END data_out[88]
  PIN data_out[89]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 2.673000 ;
    PORT
      LAYER met3 ;
        RECT 0.000 310.120 4.000 310.720 ;
    END
  END data_out[89]
  PIN data_out[8]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 2.673000 ;
    PORT
      LAYER met3 ;
        RECT 0.000 89.800 4.000 90.400 ;
    END
  END data_out[8]
  PIN data_out[90]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 2.673000 ;
    PORT
      LAYER met3 ;
        RECT 0.000 312.840 4.000 313.440 ;
    END
  END data_out[90]
  PIN data_out[91]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 2.673000 ;
    PORT
      LAYER met3 ;
        RECT 0.000 315.560 4.000 316.160 ;
    END
  END data_out[91]
  PIN data_out[92]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 2.673000 ;
    PORT
      LAYER met3 ;
        RECT 0.000 318.280 4.000 318.880 ;
    END
  END data_out[92]
  PIN data_out[93]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 2.673000 ;
    PORT
      LAYER met3 ;
        RECT 0.000 321.000 4.000 321.600 ;
    END
  END data_out[93]
  PIN data_out[94]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 2.673000 ;
    PORT
      LAYER met3 ;
        RECT 0.000 323.720 4.000 324.320 ;
    END
  END data_out[94]
  PIN data_out[95]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 2.673000 ;
    PORT
      LAYER met3 ;
        RECT 0.000 326.440 4.000 327.040 ;
    END
  END data_out[95]
  PIN data_out[96]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 2.673000 ;
    PORT
      LAYER met3 ;
        RECT 0.000 329.160 4.000 329.760 ;
    END
  END data_out[96]
  PIN data_out[97]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 2.673000 ;
    PORT
      LAYER met3 ;
        RECT 0.000 331.880 4.000 332.480 ;
    END
  END data_out[97]
  PIN data_out[98]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 2.673000 ;
    PORT
      LAYER met3 ;
        RECT 0.000 334.600 4.000 335.200 ;
    END
  END data_out[98]
  PIN data_out[99]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 2.673000 ;
    PORT
      LAYER met3 ;
        RECT 0.000 337.320 4.000 337.920 ;
    END
  END data_out[99]
  PIN data_out[9]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 2.673000 ;
    PORT
      LAYER met3 ;
        RECT 0.000 92.520 4.000 93.120 ;
    END
  END data_out[9]
  PIN done
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 2.673000 ;
    PORT
      LAYER met2 ;
        RECT 433.870 585.870 434.150 589.870 ;
    END
  END done
  PIN enable
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.126000 ;
    ANTENNADIFFAREA 0.434700 ;
    PORT
      LAYER met2 ;
        RECT 241.130 0.000 241.410 4.000 ;
    END
  END enable
  PIN ki
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.126000 ;
    ANTENNADIFFAREA 0.434700 ;
    PORT
      LAYER met2 ;
        RECT 529.550 0.000 529.830 4.000 ;
    END
  END ki
  PIN load_data
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.126000 ;
    ANTENNADIFFAREA 0.434700 ;
    PORT
      LAYER met2 ;
        RECT 337.270 0.000 337.550 4.000 ;
    END
  END load_data
  PIN load_status[0]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.126000 ;
    ANTENNADIFFAREA 0.434700 ;
    PORT
      LAYER met3 ;
        RECT 575.150 512.760 579.150 513.360 ;
    END
  END load_status[0]
  PIN load_status[1]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.126000 ;
    ANTENNADIFFAREA 0.434700 ;
    PORT
      LAYER met3 ;
        RECT 575.150 515.480 579.150 516.080 ;
    END
  END load_status[1]
  PIN load_status[2]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.126000 ;
    ANTENNADIFFAREA 0.434700 ;
    PORT
      LAYER met3 ;
        RECT 575.150 518.200 579.150 518.800 ;
    END
  END load_status[2]
  PIN next_key
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 2.673000 ;
    PORT
      LAYER met2 ;
        RECT 144.530 585.870 144.810 589.870 ;
    END
  END next_key
  PIN rst
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.196500 ;
    ANTENNADIFFAREA 0.434700 ;
    PORT
      LAYER met2 ;
        RECT 144.990 0.000 145.270 4.000 ;
    END
  END rst
  PIN trigLoad
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.126000 ;
    ANTENNADIFFAREA 0.434700 ;
    PORT
      LAYER met2 ;
        RECT 433.410 0.000 433.690 4.000 ;
    END
  END trigLoad
  PIN vccd2
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER met4 ;
        RECT 21.040 10.640 22.640 576.880 ;
    END
    PORT
      LAYER met4 ;
        RECT 174.640 10.640 176.240 576.880 ;
    END
    PORT
      LAYER met4 ;
        RECT 328.240 10.640 329.840 576.880 ;
    END
    PORT
      LAYER met4 ;
        RECT 481.840 10.640 483.440 576.880 ;
    END
  END vccd2
  PIN vssd2
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER met4 ;
        RECT 97.840 10.640 99.440 576.880 ;
    END
    PORT
      LAYER met4 ;
        RECT 251.440 10.640 253.040 576.880 ;
    END
    PORT
      LAYER met4 ;
        RECT 405.040 10.640 406.640 576.880 ;
    END
    PORT
      LAYER met4 ;
        RECT 558.640 10.640 560.240 576.880 ;
    END
  END vssd2
  OBS
      LAYER li1 ;
        RECT 5.520 10.795 573.620 576.725 ;
      LAYER met1 ;
        RECT 5.520 10.640 579.070 578.980 ;
      LAYER met2 ;
        RECT 6.070 585.590 144.250 585.870 ;
        RECT 145.090 585.590 433.590 585.870 ;
        RECT 434.430 585.590 579.050 585.870 ;
        RECT 6.070 4.280 579.050 585.590 ;
        RECT 6.070 3.670 48.570 4.280 ;
        RECT 49.410 3.670 144.710 4.280 ;
        RECT 145.550 3.670 240.850 4.280 ;
        RECT 241.690 3.670 336.990 4.280 ;
        RECT 337.830 3.670 433.130 4.280 ;
        RECT 433.970 3.670 529.270 4.280 ;
        RECT 530.110 3.670 579.050 4.280 ;
      LAYER met3 ;
        RECT 4.000 520.560 579.075 576.805 ;
        RECT 4.400 519.200 579.075 520.560 ;
        RECT 4.400 519.160 574.750 519.200 ;
        RECT 4.000 517.840 574.750 519.160 ;
        RECT 4.400 517.800 574.750 517.840 ;
        RECT 4.400 516.480 579.075 517.800 ;
        RECT 4.400 516.440 574.750 516.480 ;
        RECT 4.000 515.120 574.750 516.440 ;
        RECT 4.400 515.080 574.750 515.120 ;
        RECT 4.400 513.760 579.075 515.080 ;
        RECT 4.400 513.720 574.750 513.760 ;
        RECT 4.000 512.400 574.750 513.720 ;
        RECT 4.400 512.360 574.750 512.400 ;
        RECT 4.400 511.040 579.075 512.360 ;
        RECT 4.400 511.000 574.750 511.040 ;
        RECT 4.000 509.680 574.750 511.000 ;
        RECT 4.400 509.640 574.750 509.680 ;
        RECT 4.400 508.320 579.075 509.640 ;
        RECT 4.400 508.280 574.750 508.320 ;
        RECT 4.000 506.960 574.750 508.280 ;
        RECT 4.400 506.920 574.750 506.960 ;
        RECT 4.400 505.600 579.075 506.920 ;
        RECT 4.400 505.560 574.750 505.600 ;
        RECT 4.000 504.240 574.750 505.560 ;
        RECT 4.400 504.200 574.750 504.240 ;
        RECT 4.400 502.880 579.075 504.200 ;
        RECT 4.400 502.840 574.750 502.880 ;
        RECT 4.000 501.520 574.750 502.840 ;
        RECT 4.400 501.480 574.750 501.520 ;
        RECT 4.400 500.160 579.075 501.480 ;
        RECT 4.400 500.120 574.750 500.160 ;
        RECT 4.000 498.800 574.750 500.120 ;
        RECT 4.400 498.760 574.750 498.800 ;
        RECT 4.400 497.440 579.075 498.760 ;
        RECT 4.400 497.400 574.750 497.440 ;
        RECT 4.000 496.080 574.750 497.400 ;
        RECT 4.400 496.040 574.750 496.080 ;
        RECT 4.400 494.720 579.075 496.040 ;
        RECT 4.400 494.680 574.750 494.720 ;
        RECT 4.000 493.360 574.750 494.680 ;
        RECT 4.400 493.320 574.750 493.360 ;
        RECT 4.400 492.000 579.075 493.320 ;
        RECT 4.400 491.960 574.750 492.000 ;
        RECT 4.000 490.640 574.750 491.960 ;
        RECT 4.400 490.600 574.750 490.640 ;
        RECT 4.400 489.280 579.075 490.600 ;
        RECT 4.400 489.240 574.750 489.280 ;
        RECT 4.000 487.920 574.750 489.240 ;
        RECT 4.400 487.880 574.750 487.920 ;
        RECT 4.400 486.560 579.075 487.880 ;
        RECT 4.400 486.520 574.750 486.560 ;
        RECT 4.000 485.200 574.750 486.520 ;
        RECT 4.400 485.160 574.750 485.200 ;
        RECT 4.400 483.840 579.075 485.160 ;
        RECT 4.400 483.800 574.750 483.840 ;
        RECT 4.000 482.480 574.750 483.800 ;
        RECT 4.400 482.440 574.750 482.480 ;
        RECT 4.400 481.120 579.075 482.440 ;
        RECT 4.400 481.080 574.750 481.120 ;
        RECT 4.000 479.760 574.750 481.080 ;
        RECT 4.400 479.720 574.750 479.760 ;
        RECT 4.400 478.400 579.075 479.720 ;
        RECT 4.400 478.360 574.750 478.400 ;
        RECT 4.000 477.040 574.750 478.360 ;
        RECT 4.400 477.000 574.750 477.040 ;
        RECT 4.400 475.680 579.075 477.000 ;
        RECT 4.400 475.640 574.750 475.680 ;
        RECT 4.000 474.320 574.750 475.640 ;
        RECT 4.400 474.280 574.750 474.320 ;
        RECT 4.400 472.960 579.075 474.280 ;
        RECT 4.400 472.920 574.750 472.960 ;
        RECT 4.000 471.600 574.750 472.920 ;
        RECT 4.400 471.560 574.750 471.600 ;
        RECT 4.400 470.240 579.075 471.560 ;
        RECT 4.400 470.200 574.750 470.240 ;
        RECT 4.000 468.880 574.750 470.200 ;
        RECT 4.400 468.840 574.750 468.880 ;
        RECT 4.400 467.520 579.075 468.840 ;
        RECT 4.400 467.480 574.750 467.520 ;
        RECT 4.000 466.160 574.750 467.480 ;
        RECT 4.400 466.120 574.750 466.160 ;
        RECT 4.400 464.800 579.075 466.120 ;
        RECT 4.400 464.760 574.750 464.800 ;
        RECT 4.000 463.440 574.750 464.760 ;
        RECT 4.400 463.400 574.750 463.440 ;
        RECT 4.400 462.080 579.075 463.400 ;
        RECT 4.400 462.040 574.750 462.080 ;
        RECT 4.000 460.720 574.750 462.040 ;
        RECT 4.400 460.680 574.750 460.720 ;
        RECT 4.400 459.360 579.075 460.680 ;
        RECT 4.400 459.320 574.750 459.360 ;
        RECT 4.000 458.000 574.750 459.320 ;
        RECT 4.400 457.960 574.750 458.000 ;
        RECT 4.400 456.640 579.075 457.960 ;
        RECT 4.400 456.600 574.750 456.640 ;
        RECT 4.000 455.280 574.750 456.600 ;
        RECT 4.400 455.240 574.750 455.280 ;
        RECT 4.400 453.920 579.075 455.240 ;
        RECT 4.400 453.880 574.750 453.920 ;
        RECT 4.000 452.560 574.750 453.880 ;
        RECT 4.400 452.520 574.750 452.560 ;
        RECT 4.400 451.200 579.075 452.520 ;
        RECT 4.400 451.160 574.750 451.200 ;
        RECT 4.000 449.840 574.750 451.160 ;
        RECT 4.400 449.800 574.750 449.840 ;
        RECT 4.400 448.480 579.075 449.800 ;
        RECT 4.400 448.440 574.750 448.480 ;
        RECT 4.000 447.120 574.750 448.440 ;
        RECT 4.400 447.080 574.750 447.120 ;
        RECT 4.400 445.760 579.075 447.080 ;
        RECT 4.400 445.720 574.750 445.760 ;
        RECT 4.000 444.400 574.750 445.720 ;
        RECT 4.400 444.360 574.750 444.400 ;
        RECT 4.400 443.040 579.075 444.360 ;
        RECT 4.400 443.000 574.750 443.040 ;
        RECT 4.000 441.680 574.750 443.000 ;
        RECT 4.400 441.640 574.750 441.680 ;
        RECT 4.400 440.320 579.075 441.640 ;
        RECT 4.400 440.280 574.750 440.320 ;
        RECT 4.000 438.960 574.750 440.280 ;
        RECT 4.400 438.920 574.750 438.960 ;
        RECT 4.400 437.600 579.075 438.920 ;
        RECT 4.400 437.560 574.750 437.600 ;
        RECT 4.000 436.240 574.750 437.560 ;
        RECT 4.400 436.200 574.750 436.240 ;
        RECT 4.400 434.880 579.075 436.200 ;
        RECT 4.400 434.840 574.750 434.880 ;
        RECT 4.000 433.520 574.750 434.840 ;
        RECT 4.400 433.480 574.750 433.520 ;
        RECT 4.400 432.160 579.075 433.480 ;
        RECT 4.400 432.120 574.750 432.160 ;
        RECT 4.000 430.800 574.750 432.120 ;
        RECT 4.400 430.760 574.750 430.800 ;
        RECT 4.400 429.440 579.075 430.760 ;
        RECT 4.400 429.400 574.750 429.440 ;
        RECT 4.000 428.080 574.750 429.400 ;
        RECT 4.400 428.040 574.750 428.080 ;
        RECT 4.400 426.720 579.075 428.040 ;
        RECT 4.400 426.680 574.750 426.720 ;
        RECT 4.000 425.360 574.750 426.680 ;
        RECT 4.400 425.320 574.750 425.360 ;
        RECT 4.400 424.000 579.075 425.320 ;
        RECT 4.400 423.960 574.750 424.000 ;
        RECT 4.000 422.640 574.750 423.960 ;
        RECT 4.400 422.600 574.750 422.640 ;
        RECT 4.400 421.280 579.075 422.600 ;
        RECT 4.400 421.240 574.750 421.280 ;
        RECT 4.000 419.920 574.750 421.240 ;
        RECT 4.400 419.880 574.750 419.920 ;
        RECT 4.400 418.560 579.075 419.880 ;
        RECT 4.400 418.520 574.750 418.560 ;
        RECT 4.000 417.200 574.750 418.520 ;
        RECT 4.400 417.160 574.750 417.200 ;
        RECT 4.400 415.840 579.075 417.160 ;
        RECT 4.400 415.800 574.750 415.840 ;
        RECT 4.000 414.480 574.750 415.800 ;
        RECT 4.400 414.440 574.750 414.480 ;
        RECT 4.400 413.120 579.075 414.440 ;
        RECT 4.400 413.080 574.750 413.120 ;
        RECT 4.000 411.760 574.750 413.080 ;
        RECT 4.400 411.720 574.750 411.760 ;
        RECT 4.400 410.400 579.075 411.720 ;
        RECT 4.400 410.360 574.750 410.400 ;
        RECT 4.000 409.040 574.750 410.360 ;
        RECT 4.400 409.000 574.750 409.040 ;
        RECT 4.400 407.680 579.075 409.000 ;
        RECT 4.400 407.640 574.750 407.680 ;
        RECT 4.000 406.320 574.750 407.640 ;
        RECT 4.400 406.280 574.750 406.320 ;
        RECT 4.400 404.960 579.075 406.280 ;
        RECT 4.400 404.920 574.750 404.960 ;
        RECT 4.000 403.600 574.750 404.920 ;
        RECT 4.400 403.560 574.750 403.600 ;
        RECT 4.400 402.240 579.075 403.560 ;
        RECT 4.400 402.200 574.750 402.240 ;
        RECT 4.000 400.880 574.750 402.200 ;
        RECT 4.400 400.840 574.750 400.880 ;
        RECT 4.400 399.520 579.075 400.840 ;
        RECT 4.400 399.480 574.750 399.520 ;
        RECT 4.000 398.160 574.750 399.480 ;
        RECT 4.400 398.120 574.750 398.160 ;
        RECT 4.400 396.800 579.075 398.120 ;
        RECT 4.400 396.760 574.750 396.800 ;
        RECT 4.000 395.440 574.750 396.760 ;
        RECT 4.400 395.400 574.750 395.440 ;
        RECT 4.400 394.080 579.075 395.400 ;
        RECT 4.400 394.040 574.750 394.080 ;
        RECT 4.000 392.720 574.750 394.040 ;
        RECT 4.400 392.680 574.750 392.720 ;
        RECT 4.400 391.360 579.075 392.680 ;
        RECT 4.400 391.320 574.750 391.360 ;
        RECT 4.000 390.000 574.750 391.320 ;
        RECT 4.400 389.960 574.750 390.000 ;
        RECT 4.400 388.640 579.075 389.960 ;
        RECT 4.400 388.600 574.750 388.640 ;
        RECT 4.000 387.280 574.750 388.600 ;
        RECT 4.400 387.240 574.750 387.280 ;
        RECT 4.400 385.920 579.075 387.240 ;
        RECT 4.400 385.880 574.750 385.920 ;
        RECT 4.000 384.560 574.750 385.880 ;
        RECT 4.400 384.520 574.750 384.560 ;
        RECT 4.400 383.200 579.075 384.520 ;
        RECT 4.400 383.160 574.750 383.200 ;
        RECT 4.000 381.840 574.750 383.160 ;
        RECT 4.400 381.800 574.750 381.840 ;
        RECT 4.400 380.480 579.075 381.800 ;
        RECT 4.400 380.440 574.750 380.480 ;
        RECT 4.000 379.120 574.750 380.440 ;
        RECT 4.400 379.080 574.750 379.120 ;
        RECT 4.400 377.760 579.075 379.080 ;
        RECT 4.400 377.720 574.750 377.760 ;
        RECT 4.000 376.400 574.750 377.720 ;
        RECT 4.400 376.360 574.750 376.400 ;
        RECT 4.400 375.040 579.075 376.360 ;
        RECT 4.400 375.000 574.750 375.040 ;
        RECT 4.000 373.680 574.750 375.000 ;
        RECT 4.400 373.640 574.750 373.680 ;
        RECT 4.400 372.320 579.075 373.640 ;
        RECT 4.400 372.280 574.750 372.320 ;
        RECT 4.000 370.960 574.750 372.280 ;
        RECT 4.400 370.920 574.750 370.960 ;
        RECT 4.400 369.600 579.075 370.920 ;
        RECT 4.400 369.560 574.750 369.600 ;
        RECT 4.000 368.240 574.750 369.560 ;
        RECT 4.400 368.200 574.750 368.240 ;
        RECT 4.400 366.880 579.075 368.200 ;
        RECT 4.400 366.840 574.750 366.880 ;
        RECT 4.000 365.520 574.750 366.840 ;
        RECT 4.400 365.480 574.750 365.520 ;
        RECT 4.400 364.160 579.075 365.480 ;
        RECT 4.400 364.120 574.750 364.160 ;
        RECT 4.000 362.800 574.750 364.120 ;
        RECT 4.400 362.760 574.750 362.800 ;
        RECT 4.400 361.440 579.075 362.760 ;
        RECT 4.400 361.400 574.750 361.440 ;
        RECT 4.000 360.080 574.750 361.400 ;
        RECT 4.400 360.040 574.750 360.080 ;
        RECT 4.400 358.720 579.075 360.040 ;
        RECT 4.400 358.680 574.750 358.720 ;
        RECT 4.000 357.360 574.750 358.680 ;
        RECT 4.400 357.320 574.750 357.360 ;
        RECT 4.400 356.000 579.075 357.320 ;
        RECT 4.400 355.960 574.750 356.000 ;
        RECT 4.000 354.640 574.750 355.960 ;
        RECT 4.400 354.600 574.750 354.640 ;
        RECT 4.400 353.280 579.075 354.600 ;
        RECT 4.400 353.240 574.750 353.280 ;
        RECT 4.000 351.920 574.750 353.240 ;
        RECT 4.400 351.880 574.750 351.920 ;
        RECT 4.400 350.560 579.075 351.880 ;
        RECT 4.400 350.520 574.750 350.560 ;
        RECT 4.000 349.200 574.750 350.520 ;
        RECT 4.400 349.160 574.750 349.200 ;
        RECT 4.400 347.840 579.075 349.160 ;
        RECT 4.400 347.800 574.750 347.840 ;
        RECT 4.000 346.480 574.750 347.800 ;
        RECT 4.400 346.440 574.750 346.480 ;
        RECT 4.400 345.120 579.075 346.440 ;
        RECT 4.400 345.080 574.750 345.120 ;
        RECT 4.000 343.760 574.750 345.080 ;
        RECT 4.400 343.720 574.750 343.760 ;
        RECT 4.400 342.400 579.075 343.720 ;
        RECT 4.400 342.360 574.750 342.400 ;
        RECT 4.000 341.040 574.750 342.360 ;
        RECT 4.400 341.000 574.750 341.040 ;
        RECT 4.400 339.680 579.075 341.000 ;
        RECT 4.400 339.640 574.750 339.680 ;
        RECT 4.000 338.320 574.750 339.640 ;
        RECT 4.400 338.280 574.750 338.320 ;
        RECT 4.400 336.960 579.075 338.280 ;
        RECT 4.400 336.920 574.750 336.960 ;
        RECT 4.000 335.600 574.750 336.920 ;
        RECT 4.400 335.560 574.750 335.600 ;
        RECT 4.400 334.240 579.075 335.560 ;
        RECT 4.400 334.200 574.750 334.240 ;
        RECT 4.000 332.880 574.750 334.200 ;
        RECT 4.400 332.840 574.750 332.880 ;
        RECT 4.400 331.520 579.075 332.840 ;
        RECT 4.400 331.480 574.750 331.520 ;
        RECT 4.000 330.160 574.750 331.480 ;
        RECT 4.400 330.120 574.750 330.160 ;
        RECT 4.400 328.800 579.075 330.120 ;
        RECT 4.400 328.760 574.750 328.800 ;
        RECT 4.000 327.440 574.750 328.760 ;
        RECT 4.400 327.400 574.750 327.440 ;
        RECT 4.400 326.080 579.075 327.400 ;
        RECT 4.400 326.040 574.750 326.080 ;
        RECT 4.000 324.720 574.750 326.040 ;
        RECT 4.400 324.680 574.750 324.720 ;
        RECT 4.400 323.360 579.075 324.680 ;
        RECT 4.400 323.320 574.750 323.360 ;
        RECT 4.000 322.000 574.750 323.320 ;
        RECT 4.400 321.960 574.750 322.000 ;
        RECT 4.400 320.640 579.075 321.960 ;
        RECT 4.400 320.600 574.750 320.640 ;
        RECT 4.000 319.280 574.750 320.600 ;
        RECT 4.400 319.240 574.750 319.280 ;
        RECT 4.400 317.920 579.075 319.240 ;
        RECT 4.400 317.880 574.750 317.920 ;
        RECT 4.000 316.560 574.750 317.880 ;
        RECT 4.400 316.520 574.750 316.560 ;
        RECT 4.400 315.200 579.075 316.520 ;
        RECT 4.400 315.160 574.750 315.200 ;
        RECT 4.000 313.840 574.750 315.160 ;
        RECT 4.400 313.800 574.750 313.840 ;
        RECT 4.400 312.480 579.075 313.800 ;
        RECT 4.400 312.440 574.750 312.480 ;
        RECT 4.000 311.120 574.750 312.440 ;
        RECT 4.400 311.080 574.750 311.120 ;
        RECT 4.400 309.760 579.075 311.080 ;
        RECT 4.400 309.720 574.750 309.760 ;
        RECT 4.000 308.400 574.750 309.720 ;
        RECT 4.400 308.360 574.750 308.400 ;
        RECT 4.400 307.040 579.075 308.360 ;
        RECT 4.400 307.000 574.750 307.040 ;
        RECT 4.000 305.680 574.750 307.000 ;
        RECT 4.400 305.640 574.750 305.680 ;
        RECT 4.400 304.320 579.075 305.640 ;
        RECT 4.400 304.280 574.750 304.320 ;
        RECT 4.000 302.960 574.750 304.280 ;
        RECT 4.400 302.920 574.750 302.960 ;
        RECT 4.400 301.600 579.075 302.920 ;
        RECT 4.400 301.560 574.750 301.600 ;
        RECT 4.000 300.240 574.750 301.560 ;
        RECT 4.400 300.200 574.750 300.240 ;
        RECT 4.400 298.880 579.075 300.200 ;
        RECT 4.400 298.840 574.750 298.880 ;
        RECT 4.000 297.520 574.750 298.840 ;
        RECT 4.400 297.480 574.750 297.520 ;
        RECT 4.400 296.160 579.075 297.480 ;
        RECT 4.400 296.120 574.750 296.160 ;
        RECT 4.000 294.800 574.750 296.120 ;
        RECT 4.400 294.760 574.750 294.800 ;
        RECT 4.400 293.440 579.075 294.760 ;
        RECT 4.400 293.400 574.750 293.440 ;
        RECT 4.000 292.080 574.750 293.400 ;
        RECT 4.400 292.040 574.750 292.080 ;
        RECT 4.400 290.720 579.075 292.040 ;
        RECT 4.400 290.680 574.750 290.720 ;
        RECT 4.000 289.360 574.750 290.680 ;
        RECT 4.400 289.320 574.750 289.360 ;
        RECT 4.400 288.000 579.075 289.320 ;
        RECT 4.400 287.960 574.750 288.000 ;
        RECT 4.000 286.640 574.750 287.960 ;
        RECT 4.400 286.600 574.750 286.640 ;
        RECT 4.400 285.280 579.075 286.600 ;
        RECT 4.400 285.240 574.750 285.280 ;
        RECT 4.000 283.920 574.750 285.240 ;
        RECT 4.400 283.880 574.750 283.920 ;
        RECT 4.400 282.560 579.075 283.880 ;
        RECT 4.400 282.520 574.750 282.560 ;
        RECT 4.000 281.200 574.750 282.520 ;
        RECT 4.400 281.160 574.750 281.200 ;
        RECT 4.400 279.840 579.075 281.160 ;
        RECT 4.400 279.800 574.750 279.840 ;
        RECT 4.000 278.480 574.750 279.800 ;
        RECT 4.400 278.440 574.750 278.480 ;
        RECT 4.400 277.120 579.075 278.440 ;
        RECT 4.400 277.080 574.750 277.120 ;
        RECT 4.000 275.760 574.750 277.080 ;
        RECT 4.400 275.720 574.750 275.760 ;
        RECT 4.400 274.400 579.075 275.720 ;
        RECT 4.400 274.360 574.750 274.400 ;
        RECT 4.000 273.040 574.750 274.360 ;
        RECT 4.400 273.000 574.750 273.040 ;
        RECT 4.400 271.680 579.075 273.000 ;
        RECT 4.400 271.640 574.750 271.680 ;
        RECT 4.000 270.320 574.750 271.640 ;
        RECT 4.400 270.280 574.750 270.320 ;
        RECT 4.400 268.960 579.075 270.280 ;
        RECT 4.400 268.920 574.750 268.960 ;
        RECT 4.000 267.600 574.750 268.920 ;
        RECT 4.400 267.560 574.750 267.600 ;
        RECT 4.400 266.240 579.075 267.560 ;
        RECT 4.400 266.200 574.750 266.240 ;
        RECT 4.000 264.880 574.750 266.200 ;
        RECT 4.400 264.840 574.750 264.880 ;
        RECT 4.400 263.520 579.075 264.840 ;
        RECT 4.400 263.480 574.750 263.520 ;
        RECT 4.000 262.160 574.750 263.480 ;
        RECT 4.400 262.120 574.750 262.160 ;
        RECT 4.400 260.800 579.075 262.120 ;
        RECT 4.400 260.760 574.750 260.800 ;
        RECT 4.000 259.440 574.750 260.760 ;
        RECT 4.400 259.400 574.750 259.440 ;
        RECT 4.400 258.080 579.075 259.400 ;
        RECT 4.400 258.040 574.750 258.080 ;
        RECT 4.000 256.720 574.750 258.040 ;
        RECT 4.400 256.680 574.750 256.720 ;
        RECT 4.400 255.360 579.075 256.680 ;
        RECT 4.400 255.320 574.750 255.360 ;
        RECT 4.000 254.000 574.750 255.320 ;
        RECT 4.400 253.960 574.750 254.000 ;
        RECT 4.400 252.640 579.075 253.960 ;
        RECT 4.400 252.600 574.750 252.640 ;
        RECT 4.000 251.280 574.750 252.600 ;
        RECT 4.400 251.240 574.750 251.280 ;
        RECT 4.400 249.920 579.075 251.240 ;
        RECT 4.400 249.880 574.750 249.920 ;
        RECT 4.000 248.560 574.750 249.880 ;
        RECT 4.400 248.520 574.750 248.560 ;
        RECT 4.400 247.200 579.075 248.520 ;
        RECT 4.400 247.160 574.750 247.200 ;
        RECT 4.000 245.840 574.750 247.160 ;
        RECT 4.400 245.800 574.750 245.840 ;
        RECT 4.400 244.480 579.075 245.800 ;
        RECT 4.400 244.440 574.750 244.480 ;
        RECT 4.000 243.120 574.750 244.440 ;
        RECT 4.400 243.080 574.750 243.120 ;
        RECT 4.400 241.760 579.075 243.080 ;
        RECT 4.400 241.720 574.750 241.760 ;
        RECT 4.000 240.400 574.750 241.720 ;
        RECT 4.400 240.360 574.750 240.400 ;
        RECT 4.400 239.040 579.075 240.360 ;
        RECT 4.400 239.000 574.750 239.040 ;
        RECT 4.000 237.680 574.750 239.000 ;
        RECT 4.400 237.640 574.750 237.680 ;
        RECT 4.400 236.320 579.075 237.640 ;
        RECT 4.400 236.280 574.750 236.320 ;
        RECT 4.000 234.960 574.750 236.280 ;
        RECT 4.400 234.920 574.750 234.960 ;
        RECT 4.400 233.600 579.075 234.920 ;
        RECT 4.400 233.560 574.750 233.600 ;
        RECT 4.000 232.240 574.750 233.560 ;
        RECT 4.400 232.200 574.750 232.240 ;
        RECT 4.400 230.880 579.075 232.200 ;
        RECT 4.400 230.840 574.750 230.880 ;
        RECT 4.000 229.520 574.750 230.840 ;
        RECT 4.400 229.480 574.750 229.520 ;
        RECT 4.400 228.160 579.075 229.480 ;
        RECT 4.400 228.120 574.750 228.160 ;
        RECT 4.000 226.800 574.750 228.120 ;
        RECT 4.400 226.760 574.750 226.800 ;
        RECT 4.400 225.440 579.075 226.760 ;
        RECT 4.400 225.400 574.750 225.440 ;
        RECT 4.000 224.080 574.750 225.400 ;
        RECT 4.400 224.040 574.750 224.080 ;
        RECT 4.400 222.720 579.075 224.040 ;
        RECT 4.400 222.680 574.750 222.720 ;
        RECT 4.000 221.360 574.750 222.680 ;
        RECT 4.400 221.320 574.750 221.360 ;
        RECT 4.400 220.000 579.075 221.320 ;
        RECT 4.400 219.960 574.750 220.000 ;
        RECT 4.000 218.640 574.750 219.960 ;
        RECT 4.400 218.600 574.750 218.640 ;
        RECT 4.400 217.280 579.075 218.600 ;
        RECT 4.400 217.240 574.750 217.280 ;
        RECT 4.000 215.920 574.750 217.240 ;
        RECT 4.400 215.880 574.750 215.920 ;
        RECT 4.400 214.560 579.075 215.880 ;
        RECT 4.400 214.520 574.750 214.560 ;
        RECT 4.000 213.200 574.750 214.520 ;
        RECT 4.400 213.160 574.750 213.200 ;
        RECT 4.400 211.840 579.075 213.160 ;
        RECT 4.400 211.800 574.750 211.840 ;
        RECT 4.000 210.480 574.750 211.800 ;
        RECT 4.400 210.440 574.750 210.480 ;
        RECT 4.400 209.120 579.075 210.440 ;
        RECT 4.400 209.080 574.750 209.120 ;
        RECT 4.000 207.760 574.750 209.080 ;
        RECT 4.400 207.720 574.750 207.760 ;
        RECT 4.400 206.400 579.075 207.720 ;
        RECT 4.400 206.360 574.750 206.400 ;
        RECT 4.000 205.040 574.750 206.360 ;
        RECT 4.400 205.000 574.750 205.040 ;
        RECT 4.400 203.680 579.075 205.000 ;
        RECT 4.400 203.640 574.750 203.680 ;
        RECT 4.000 202.320 574.750 203.640 ;
        RECT 4.400 202.280 574.750 202.320 ;
        RECT 4.400 200.960 579.075 202.280 ;
        RECT 4.400 200.920 574.750 200.960 ;
        RECT 4.000 199.600 574.750 200.920 ;
        RECT 4.400 199.560 574.750 199.600 ;
        RECT 4.400 198.240 579.075 199.560 ;
        RECT 4.400 198.200 574.750 198.240 ;
        RECT 4.000 196.880 574.750 198.200 ;
        RECT 4.400 196.840 574.750 196.880 ;
        RECT 4.400 195.520 579.075 196.840 ;
        RECT 4.400 195.480 574.750 195.520 ;
        RECT 4.000 194.160 574.750 195.480 ;
        RECT 4.400 194.120 574.750 194.160 ;
        RECT 4.400 192.800 579.075 194.120 ;
        RECT 4.400 192.760 574.750 192.800 ;
        RECT 4.000 191.440 574.750 192.760 ;
        RECT 4.400 191.400 574.750 191.440 ;
        RECT 4.400 190.080 579.075 191.400 ;
        RECT 4.400 190.040 574.750 190.080 ;
        RECT 4.000 188.720 574.750 190.040 ;
        RECT 4.400 188.680 574.750 188.720 ;
        RECT 4.400 187.360 579.075 188.680 ;
        RECT 4.400 187.320 574.750 187.360 ;
        RECT 4.000 186.000 574.750 187.320 ;
        RECT 4.400 185.960 574.750 186.000 ;
        RECT 4.400 184.640 579.075 185.960 ;
        RECT 4.400 184.600 574.750 184.640 ;
        RECT 4.000 183.280 574.750 184.600 ;
        RECT 4.400 183.240 574.750 183.280 ;
        RECT 4.400 181.920 579.075 183.240 ;
        RECT 4.400 181.880 574.750 181.920 ;
        RECT 4.000 180.560 574.750 181.880 ;
        RECT 4.400 180.520 574.750 180.560 ;
        RECT 4.400 179.200 579.075 180.520 ;
        RECT 4.400 179.160 574.750 179.200 ;
        RECT 4.000 177.840 574.750 179.160 ;
        RECT 4.400 177.800 574.750 177.840 ;
        RECT 4.400 176.480 579.075 177.800 ;
        RECT 4.400 176.440 574.750 176.480 ;
        RECT 4.000 175.120 574.750 176.440 ;
        RECT 4.400 175.080 574.750 175.120 ;
        RECT 4.400 173.760 579.075 175.080 ;
        RECT 4.400 173.720 574.750 173.760 ;
        RECT 4.000 172.400 574.750 173.720 ;
        RECT 4.400 172.360 574.750 172.400 ;
        RECT 4.400 171.040 579.075 172.360 ;
        RECT 4.400 171.000 574.750 171.040 ;
        RECT 4.000 169.680 574.750 171.000 ;
        RECT 4.400 169.640 574.750 169.680 ;
        RECT 4.400 168.320 579.075 169.640 ;
        RECT 4.400 168.280 574.750 168.320 ;
        RECT 4.000 166.960 574.750 168.280 ;
        RECT 4.400 166.920 574.750 166.960 ;
        RECT 4.400 165.600 579.075 166.920 ;
        RECT 4.400 165.560 574.750 165.600 ;
        RECT 4.000 164.240 574.750 165.560 ;
        RECT 4.400 164.200 574.750 164.240 ;
        RECT 4.400 162.880 579.075 164.200 ;
        RECT 4.400 162.840 574.750 162.880 ;
        RECT 4.000 161.520 574.750 162.840 ;
        RECT 4.400 161.480 574.750 161.520 ;
        RECT 4.400 160.160 579.075 161.480 ;
        RECT 4.400 160.120 574.750 160.160 ;
        RECT 4.000 158.800 574.750 160.120 ;
        RECT 4.400 158.760 574.750 158.800 ;
        RECT 4.400 157.440 579.075 158.760 ;
        RECT 4.400 157.400 574.750 157.440 ;
        RECT 4.000 156.080 574.750 157.400 ;
        RECT 4.400 156.040 574.750 156.080 ;
        RECT 4.400 154.720 579.075 156.040 ;
        RECT 4.400 154.680 574.750 154.720 ;
        RECT 4.000 153.360 574.750 154.680 ;
        RECT 4.400 153.320 574.750 153.360 ;
        RECT 4.400 152.000 579.075 153.320 ;
        RECT 4.400 151.960 574.750 152.000 ;
        RECT 4.000 150.640 574.750 151.960 ;
        RECT 4.400 150.600 574.750 150.640 ;
        RECT 4.400 149.280 579.075 150.600 ;
        RECT 4.400 149.240 574.750 149.280 ;
        RECT 4.000 147.920 574.750 149.240 ;
        RECT 4.400 147.880 574.750 147.920 ;
        RECT 4.400 146.560 579.075 147.880 ;
        RECT 4.400 146.520 574.750 146.560 ;
        RECT 4.000 145.200 574.750 146.520 ;
        RECT 4.400 145.160 574.750 145.200 ;
        RECT 4.400 143.840 579.075 145.160 ;
        RECT 4.400 143.800 574.750 143.840 ;
        RECT 4.000 142.480 574.750 143.800 ;
        RECT 4.400 142.440 574.750 142.480 ;
        RECT 4.400 141.120 579.075 142.440 ;
        RECT 4.400 141.080 574.750 141.120 ;
        RECT 4.000 139.760 574.750 141.080 ;
        RECT 4.400 139.720 574.750 139.760 ;
        RECT 4.400 138.400 579.075 139.720 ;
        RECT 4.400 138.360 574.750 138.400 ;
        RECT 4.000 137.040 574.750 138.360 ;
        RECT 4.400 137.000 574.750 137.040 ;
        RECT 4.400 135.680 579.075 137.000 ;
        RECT 4.400 135.640 574.750 135.680 ;
        RECT 4.000 134.320 574.750 135.640 ;
        RECT 4.400 134.280 574.750 134.320 ;
        RECT 4.400 132.960 579.075 134.280 ;
        RECT 4.400 132.920 574.750 132.960 ;
        RECT 4.000 131.600 574.750 132.920 ;
        RECT 4.400 131.560 574.750 131.600 ;
        RECT 4.400 130.240 579.075 131.560 ;
        RECT 4.400 130.200 574.750 130.240 ;
        RECT 4.000 128.880 574.750 130.200 ;
        RECT 4.400 128.840 574.750 128.880 ;
        RECT 4.400 127.520 579.075 128.840 ;
        RECT 4.400 127.480 574.750 127.520 ;
        RECT 4.000 126.160 574.750 127.480 ;
        RECT 4.400 126.120 574.750 126.160 ;
        RECT 4.400 124.800 579.075 126.120 ;
        RECT 4.400 124.760 574.750 124.800 ;
        RECT 4.000 123.440 574.750 124.760 ;
        RECT 4.400 123.400 574.750 123.440 ;
        RECT 4.400 122.080 579.075 123.400 ;
        RECT 4.400 122.040 574.750 122.080 ;
        RECT 4.000 120.720 574.750 122.040 ;
        RECT 4.400 120.680 574.750 120.720 ;
        RECT 4.400 119.360 579.075 120.680 ;
        RECT 4.400 119.320 574.750 119.360 ;
        RECT 4.000 118.000 574.750 119.320 ;
        RECT 4.400 117.960 574.750 118.000 ;
        RECT 4.400 116.640 579.075 117.960 ;
        RECT 4.400 116.600 574.750 116.640 ;
        RECT 4.000 115.280 574.750 116.600 ;
        RECT 4.400 115.240 574.750 115.280 ;
        RECT 4.400 113.920 579.075 115.240 ;
        RECT 4.400 113.880 574.750 113.920 ;
        RECT 4.000 112.560 574.750 113.880 ;
        RECT 4.400 112.520 574.750 112.560 ;
        RECT 4.400 111.200 579.075 112.520 ;
        RECT 4.400 111.160 574.750 111.200 ;
        RECT 4.000 109.840 574.750 111.160 ;
        RECT 4.400 109.800 574.750 109.840 ;
        RECT 4.400 108.480 579.075 109.800 ;
        RECT 4.400 108.440 574.750 108.480 ;
        RECT 4.000 107.120 574.750 108.440 ;
        RECT 4.400 107.080 574.750 107.120 ;
        RECT 4.400 105.760 579.075 107.080 ;
        RECT 4.400 105.720 574.750 105.760 ;
        RECT 4.000 104.400 574.750 105.720 ;
        RECT 4.400 104.360 574.750 104.400 ;
        RECT 4.400 103.040 579.075 104.360 ;
        RECT 4.400 103.000 574.750 103.040 ;
        RECT 4.000 101.680 574.750 103.000 ;
        RECT 4.400 101.640 574.750 101.680 ;
        RECT 4.400 100.320 579.075 101.640 ;
        RECT 4.400 100.280 574.750 100.320 ;
        RECT 4.000 98.960 574.750 100.280 ;
        RECT 4.400 98.920 574.750 98.960 ;
        RECT 4.400 97.600 579.075 98.920 ;
        RECT 4.400 97.560 574.750 97.600 ;
        RECT 4.000 96.240 574.750 97.560 ;
        RECT 4.400 96.200 574.750 96.240 ;
        RECT 4.400 94.880 579.075 96.200 ;
        RECT 4.400 94.840 574.750 94.880 ;
        RECT 4.000 93.520 574.750 94.840 ;
        RECT 4.400 93.480 574.750 93.520 ;
        RECT 4.400 92.160 579.075 93.480 ;
        RECT 4.400 92.120 574.750 92.160 ;
        RECT 4.000 90.800 574.750 92.120 ;
        RECT 4.400 90.760 574.750 90.800 ;
        RECT 4.400 89.440 579.075 90.760 ;
        RECT 4.400 89.400 574.750 89.440 ;
        RECT 4.000 88.080 574.750 89.400 ;
        RECT 4.400 88.040 574.750 88.080 ;
        RECT 4.400 86.720 579.075 88.040 ;
        RECT 4.400 86.680 574.750 86.720 ;
        RECT 4.000 85.360 574.750 86.680 ;
        RECT 4.400 85.320 574.750 85.360 ;
        RECT 4.400 84.000 579.075 85.320 ;
        RECT 4.400 83.960 574.750 84.000 ;
        RECT 4.000 82.640 574.750 83.960 ;
        RECT 4.400 82.600 574.750 82.640 ;
        RECT 4.400 81.280 579.075 82.600 ;
        RECT 4.400 81.240 574.750 81.280 ;
        RECT 4.000 79.920 574.750 81.240 ;
        RECT 4.400 79.880 574.750 79.920 ;
        RECT 4.400 78.560 579.075 79.880 ;
        RECT 4.400 78.520 574.750 78.560 ;
        RECT 4.000 77.200 574.750 78.520 ;
        RECT 4.400 77.160 574.750 77.200 ;
        RECT 4.400 75.840 579.075 77.160 ;
        RECT 4.400 75.800 574.750 75.840 ;
        RECT 4.000 74.480 574.750 75.800 ;
        RECT 4.400 74.440 574.750 74.480 ;
        RECT 4.400 73.120 579.075 74.440 ;
        RECT 4.400 73.080 574.750 73.120 ;
        RECT 4.000 71.760 574.750 73.080 ;
        RECT 4.400 71.720 574.750 71.760 ;
        RECT 4.400 70.400 579.075 71.720 ;
        RECT 4.400 70.360 574.750 70.400 ;
        RECT 4.000 69.040 574.750 70.360 ;
        RECT 4.400 69.000 574.750 69.040 ;
        RECT 4.400 67.640 579.075 69.000 ;
        RECT 4.000 10.715 579.075 67.640 ;
      LAYER met4 ;
        RECT 19.615 11.735 20.640 573.065 ;
        RECT 23.040 11.735 97.440 573.065 ;
        RECT 99.840 11.735 174.240 573.065 ;
        RECT 176.640 11.735 251.040 573.065 ;
        RECT 253.440 11.735 327.840 573.065 ;
        RECT 330.240 11.735 404.640 573.065 ;
        RECT 407.040 11.735 481.440 573.065 ;
        RECT 483.840 11.735 558.240 573.065 ;
        RECT 560.640 11.735 564.585 573.065 ;
  END
END sm_bec_v3
END LIBRARY

