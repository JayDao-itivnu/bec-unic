* NGSPICE file created from user_project_wrapper.ext - technology: sky130A

* Black-box entry subcircuit for sm_bec_v3 abstract view
.subckt sm_bec_v3 becStatus[0] becStatus[1] becStatus[2] becStatus[3] clk data_in[0]
+ data_in[100] data_in[101] data_in[102] data_in[103] data_in[104] data_in[105] data_in[106]
+ data_in[107] data_in[108] data_in[109] data_in[10] data_in[110] data_in[111] data_in[112]
+ data_in[113] data_in[114] data_in[115] data_in[116] data_in[117] data_in[118] data_in[119]
+ data_in[11] data_in[120] data_in[121] data_in[122] data_in[123] data_in[124] data_in[125]
+ data_in[126] data_in[127] data_in[128] data_in[129] data_in[12] data_in[130] data_in[131]
+ data_in[132] data_in[133] data_in[134] data_in[135] data_in[136] data_in[137] data_in[138]
+ data_in[139] data_in[13] data_in[140] data_in[141] data_in[142] data_in[143] data_in[144]
+ data_in[145] data_in[146] data_in[147] data_in[148] data_in[149] data_in[14] data_in[150]
+ data_in[151] data_in[152] data_in[153] data_in[154] data_in[155] data_in[156] data_in[157]
+ data_in[158] data_in[159] data_in[15] data_in[160] data_in[161] data_in[162] data_in[16]
+ data_in[17] data_in[18] data_in[19] data_in[1] data_in[20] data_in[21] data_in[22]
+ data_in[23] data_in[24] data_in[25] data_in[26] data_in[27] data_in[28] data_in[29]
+ data_in[2] data_in[30] data_in[31] data_in[32] data_in[33] data_in[34] data_in[35]
+ data_in[36] data_in[37] data_in[38] data_in[39] data_in[3] data_in[40] data_in[41]
+ data_in[42] data_in[43] data_in[44] data_in[45] data_in[46] data_in[47] data_in[48]
+ data_in[49] data_in[4] data_in[50] data_in[51] data_in[52] data_in[53] data_in[54]
+ data_in[55] data_in[56] data_in[57] data_in[58] data_in[59] data_in[5] data_in[60]
+ data_in[61] data_in[62] data_in[63] data_in[64] data_in[65] data_in[66] data_in[67]
+ data_in[68] data_in[69] data_in[6] data_in[70] data_in[71] data_in[72] data_in[73]
+ data_in[74] data_in[75] data_in[76] data_in[77] data_in[78] data_in[79] data_in[7]
+ data_in[80] data_in[81] data_in[82] data_in[83] data_in[84] data_in[85] data_in[86]
+ data_in[87] data_in[88] data_in[89] data_in[8] data_in[90] data_in[91] data_in[92]
+ data_in[93] data_in[94] data_in[95] data_in[96] data_in[97] data_in[98] data_in[99]
+ data_in[9] data_out[0] data_out[100] data_out[101] data_out[102] data_out[103] data_out[104]
+ data_out[105] data_out[106] data_out[107] data_out[108] data_out[109] data_out[10]
+ data_out[110] data_out[111] data_out[112] data_out[113] data_out[114] data_out[115]
+ data_out[116] data_out[117] data_out[118] data_out[119] data_out[11] data_out[120]
+ data_out[121] data_out[122] data_out[123] data_out[124] data_out[125] data_out[126]
+ data_out[127] data_out[128] data_out[129] data_out[12] data_out[130] data_out[131]
+ data_out[132] data_out[133] data_out[134] data_out[135] data_out[136] data_out[137]
+ data_out[138] data_out[139] data_out[13] data_out[140] data_out[141] data_out[142]
+ data_out[143] data_out[144] data_out[145] data_out[146] data_out[147] data_out[148]
+ data_out[149] data_out[14] data_out[150] data_out[151] data_out[152] data_out[153]
+ data_out[154] data_out[155] data_out[156] data_out[157] data_out[158] data_out[159]
+ data_out[15] data_out[160] data_out[161] data_out[162] data_out[16] data_out[17]
+ data_out[18] data_out[19] data_out[1] data_out[20] data_out[21] data_out[22] data_out[23]
+ data_out[24] data_out[25] data_out[26] data_out[27] data_out[28] data_out[29] data_out[2]
+ data_out[30] data_out[31] data_out[32] data_out[33] data_out[34] data_out[35] data_out[36]
+ data_out[37] data_out[38] data_out[39] data_out[3] data_out[40] data_out[41] data_out[42]
+ data_out[43] data_out[44] data_out[45] data_out[46] data_out[47] data_out[48] data_out[49]
+ data_out[4] data_out[50] data_out[51] data_out[52] data_out[53] data_out[54] data_out[55]
+ data_out[56] data_out[57] data_out[58] data_out[59] data_out[5] data_out[60] data_out[61]
+ data_out[62] data_out[63] data_out[64] data_out[65] data_out[66] data_out[67] data_out[68]
+ data_out[69] data_out[6] data_out[70] data_out[71] data_out[72] data_out[73] data_out[74]
+ data_out[75] data_out[76] data_out[77] data_out[78] data_out[79] data_out[7] data_out[80]
+ data_out[81] data_out[82] data_out[83] data_out[84] data_out[85] data_out[86] data_out[87]
+ data_out[88] data_out[89] data_out[8] data_out[90] data_out[91] data_out[92] data_out[93]
+ data_out[94] data_out[95] data_out[96] data_out[97] data_out[98] data_out[99] data_out[9]
+ done enable ki load_data load_status[0] load_status[1] load_status[2] next_key rst
+ trigLoad vccd2 vssd2
.ends

* Black-box entry subcircuit for controller abstract view
.subckt controller becStatus[0] becStatus[1] becStatus[2] becStatus[3] data_in[0]
+ data_in[100] data_in[101] data_in[102] data_in[103] data_in[104] data_in[105] data_in[106]
+ data_in[107] data_in[108] data_in[109] data_in[10] data_in[110] data_in[111] data_in[112]
+ data_in[113] data_in[114] data_in[115] data_in[116] data_in[117] data_in[118] data_in[119]
+ data_in[11] data_in[120] data_in[121] data_in[122] data_in[123] data_in[124] data_in[125]
+ data_in[126] data_in[127] data_in[128] data_in[129] data_in[12] data_in[130] data_in[131]
+ data_in[132] data_in[133] data_in[134] data_in[135] data_in[136] data_in[137] data_in[138]
+ data_in[139] data_in[13] data_in[140] data_in[141] data_in[142] data_in[143] data_in[144]
+ data_in[145] data_in[146] data_in[147] data_in[148] data_in[149] data_in[14] data_in[150]
+ data_in[151] data_in[152] data_in[153] data_in[154] data_in[155] data_in[156] data_in[157]
+ data_in[158] data_in[159] data_in[15] data_in[160] data_in[161] data_in[162] data_in[16]
+ data_in[17] data_in[18] data_in[19] data_in[1] data_in[20] data_in[21] data_in[22]
+ data_in[23] data_in[24] data_in[25] data_in[26] data_in[27] data_in[28] data_in[29]
+ data_in[2] data_in[30] data_in[31] data_in[32] data_in[33] data_in[34] data_in[35]
+ data_in[36] data_in[37] data_in[38] data_in[39] data_in[3] data_in[40] data_in[41]
+ data_in[42] data_in[43] data_in[44] data_in[45] data_in[46] data_in[47] data_in[48]
+ data_in[49] data_in[4] data_in[50] data_in[51] data_in[52] data_in[53] data_in[54]
+ data_in[55] data_in[56] data_in[57] data_in[58] data_in[59] data_in[5] data_in[60]
+ data_in[61] data_in[62] data_in[63] data_in[64] data_in[65] data_in[66] data_in[67]
+ data_in[68] data_in[69] data_in[6] data_in[70] data_in[71] data_in[72] data_in[73]
+ data_in[74] data_in[75] data_in[76] data_in[77] data_in[78] data_in[79] data_in[7]
+ data_in[80] data_in[81] data_in[82] data_in[83] data_in[84] data_in[85] data_in[86]
+ data_in[87] data_in[88] data_in[89] data_in[8] data_in[90] data_in[91] data_in[92]
+ data_in[93] data_in[94] data_in[95] data_in[96] data_in[97] data_in[98] data_in[99]
+ data_in[9] data_out[0] data_out[100] data_out[101] data_out[102] data_out[103] data_out[104]
+ data_out[105] data_out[106] data_out[107] data_out[108] data_out[109] data_out[10]
+ data_out[110] data_out[111] data_out[112] data_out[113] data_out[114] data_out[115]
+ data_out[116] data_out[117] data_out[118] data_out[119] data_out[11] data_out[120]
+ data_out[121] data_out[122] data_out[123] data_out[124] data_out[125] data_out[126]
+ data_out[127] data_out[128] data_out[129] data_out[12] data_out[130] data_out[131]
+ data_out[132] data_out[133] data_out[134] data_out[135] data_out[136] data_out[137]
+ data_out[138] data_out[139] data_out[13] data_out[140] data_out[141] data_out[142]
+ data_out[143] data_out[144] data_out[145] data_out[146] data_out[147] data_out[148]
+ data_out[149] data_out[14] data_out[150] data_out[151] data_out[152] data_out[153]
+ data_out[154] data_out[155] data_out[156] data_out[157] data_out[158] data_out[159]
+ data_out[15] data_out[160] data_out[161] data_out[162] data_out[16] data_out[17]
+ data_out[18] data_out[19] data_out[1] data_out[20] data_out[21] data_out[22] data_out[23]
+ data_out[24] data_out[25] data_out[26] data_out[27] data_out[28] data_out[29] data_out[2]
+ data_out[30] data_out[31] data_out[32] data_out[33] data_out[34] data_out[35] data_out[36]
+ data_out[37] data_out[38] data_out[39] data_out[3] data_out[40] data_out[41] data_out[42]
+ data_out[43] data_out[44] data_out[45] data_out[46] data_out[47] data_out[48] data_out[49]
+ data_out[4] data_out[50] data_out[51] data_out[52] data_out[53] data_out[54] data_out[55]
+ data_out[56] data_out[57] data_out[58] data_out[59] data_out[5] data_out[60] data_out[61]
+ data_out[62] data_out[63] data_out[64] data_out[65] data_out[66] data_out[67] data_out[68]
+ data_out[69] data_out[6] data_out[70] data_out[71] data_out[72] data_out[73] data_out[74]
+ data_out[75] data_out[76] data_out[77] data_out[78] data_out[79] data_out[7] data_out[80]
+ data_out[81] data_out[82] data_out[83] data_out[84] data_out[85] data_out[86] data_out[87]
+ data_out[88] data_out[89] data_out[8] data_out[90] data_out[91] data_out[92] data_out[93]
+ data_out[94] data_out[95] data_out[96] data_out[97] data_out[98] data_out[99] data_out[9]
+ ki la_data_in[0] la_data_in[100] la_data_in[101] la_data_in[102] la_data_in[103]
+ la_data_in[104] la_data_in[105] la_data_in[106] la_data_in[107] la_data_in[108]
+ la_data_in[109] la_data_in[10] la_data_in[110] la_data_in[111] la_data_in[112] la_data_in[113]
+ la_data_in[114] la_data_in[115] la_data_in[116] la_data_in[117] la_data_in[118]
+ la_data_in[119] la_data_in[11] la_data_in[120] la_data_in[121] la_data_in[122] la_data_in[123]
+ la_data_in[124] la_data_in[125] la_data_in[126] la_data_in[127] la_data_in[12] la_data_in[13]
+ la_data_in[14] la_data_in[15] la_data_in[16] la_data_in[17] la_data_in[18] la_data_in[19]
+ la_data_in[1] la_data_in[20] la_data_in[21] la_data_in[22] la_data_in[23] la_data_in[24]
+ la_data_in[25] la_data_in[26] la_data_in[27] la_data_in[28] la_data_in[29] la_data_in[2]
+ la_data_in[30] la_data_in[31] la_data_in[32] la_data_in[33] la_data_in[34] la_data_in[35]
+ la_data_in[36] la_data_in[37] la_data_in[38] la_data_in[39] la_data_in[3] la_data_in[40]
+ la_data_in[41] la_data_in[42] la_data_in[43] la_data_in[44] la_data_in[45] la_data_in[46]
+ la_data_in[47] la_data_in[48] la_data_in[49] la_data_in[4] la_data_in[50] la_data_in[51]
+ la_data_in[52] la_data_in[53] la_data_in[54] la_data_in[55] la_data_in[56] la_data_in[57]
+ la_data_in[58] la_data_in[59] la_data_in[5] la_data_in[60] la_data_in[61] la_data_in[62]
+ la_data_in[63] la_data_in[64] la_data_in[65] la_data_in[66] la_data_in[67] la_data_in[68]
+ la_data_in[69] la_data_in[6] la_data_in[70] la_data_in[71] la_data_in[72] la_data_in[73]
+ la_data_in[74] la_data_in[75] la_data_in[76] la_data_in[77] la_data_in[78] la_data_in[79]
+ la_data_in[7] la_data_in[80] la_data_in[81] la_data_in[82] la_data_in[83] la_data_in[84]
+ la_data_in[85] la_data_in[86] la_data_in[87] la_data_in[88] la_data_in[89] la_data_in[8]
+ la_data_in[90] la_data_in[91] la_data_in[92] la_data_in[93] la_data_in[94] la_data_in[95]
+ la_data_in[96] la_data_in[97] la_data_in[98] la_data_in[99] la_data_in[9] la_data_out[0]
+ la_data_out[100] la_data_out[101] la_data_out[102] la_data_out[103] la_data_out[104]
+ la_data_out[105] la_data_out[106] la_data_out[107] la_data_out[108] la_data_out[109]
+ la_data_out[10] la_data_out[110] la_data_out[111] la_data_out[112] la_data_out[113]
+ la_data_out[114] la_data_out[115] la_data_out[116] la_data_out[117] la_data_out[118]
+ la_data_out[119] la_data_out[11] la_data_out[120] la_data_out[121] la_data_out[122]
+ la_data_out[123] la_data_out[124] la_data_out[125] la_data_out[126] la_data_out[127]
+ la_data_out[12] la_data_out[13] la_data_out[14] la_data_out[15] la_data_out[16]
+ la_data_out[17] la_data_out[18] la_data_out[19] la_data_out[1] la_data_out[20] la_data_out[21]
+ la_data_out[22] la_data_out[23] la_data_out[24] la_data_out[25] la_data_out[26]
+ la_data_out[27] la_data_out[28] la_data_out[29] la_data_out[2] la_data_out[30] la_data_out[31]
+ la_data_out[32] la_data_out[33] la_data_out[34] la_data_out[35] la_data_out[36]
+ la_data_out[37] la_data_out[38] la_data_out[39] la_data_out[3] la_data_out[40] la_data_out[41]
+ la_data_out[42] la_data_out[43] la_data_out[44] la_data_out[45] la_data_out[46]
+ la_data_out[47] la_data_out[48] la_data_out[49] la_data_out[4] la_data_out[50] la_data_out[51]
+ la_data_out[52] la_data_out[53] la_data_out[54] la_data_out[55] la_data_out[56]
+ la_data_out[57] la_data_out[58] la_data_out[59] la_data_out[5] la_data_out[60] la_data_out[61]
+ la_data_out[62] la_data_out[63] la_data_out[64] la_data_out[65] la_data_out[66]
+ la_data_out[67] la_data_out[68] la_data_out[69] la_data_out[6] la_data_out[70] la_data_out[71]
+ la_data_out[72] la_data_out[73] la_data_out[74] la_data_out[75] la_data_out[76]
+ la_data_out[77] la_data_out[78] la_data_out[79] la_data_out[7] la_data_out[80] la_data_out[81]
+ la_data_out[82] la_data_out[83] la_data_out[84] la_data_out[85] la_data_out[86]
+ la_data_out[87] la_data_out[88] la_data_out[89] la_data_out[8] la_data_out[90] la_data_out[91]
+ la_data_out[92] la_data_out[93] la_data_out[94] la_data_out[95] la_data_out[96]
+ la_data_out[97] la_data_out[98] la_data_out[99] la_data_out[9] la_oenb[0] la_oenb[100]
+ la_oenb[101] la_oenb[102] la_oenb[103] la_oenb[104] la_oenb[105] la_oenb[106] la_oenb[107]
+ la_oenb[108] la_oenb[109] la_oenb[10] la_oenb[110] la_oenb[111] la_oenb[112] la_oenb[113]
+ la_oenb[114] la_oenb[115] la_oenb[116] la_oenb[117] la_oenb[118] la_oenb[119] la_oenb[11]
+ la_oenb[120] la_oenb[121] la_oenb[122] la_oenb[123] la_oenb[124] la_oenb[125] la_oenb[126]
+ la_oenb[127] la_oenb[12] la_oenb[13] la_oenb[14] la_oenb[15] la_oenb[16] la_oenb[17]
+ la_oenb[18] la_oenb[19] la_oenb[1] la_oenb[20] la_oenb[21] la_oenb[22] la_oenb[23]
+ la_oenb[24] la_oenb[25] la_oenb[26] la_oenb[27] la_oenb[28] la_oenb[29] la_oenb[2]
+ la_oenb[30] la_oenb[31] la_oenb[32] la_oenb[33] la_oenb[34] la_oenb[35] la_oenb[36]
+ la_oenb[37] la_oenb[38] la_oenb[39] la_oenb[3] la_oenb[40] la_oenb[41] la_oenb[42]
+ la_oenb[43] la_oenb[44] la_oenb[45] la_oenb[46] la_oenb[47] la_oenb[48] la_oenb[49]
+ la_oenb[4] la_oenb[50] la_oenb[51] la_oenb[52] la_oenb[53] la_oenb[54] la_oenb[55]
+ la_oenb[56] la_oenb[57] la_oenb[58] la_oenb[59] la_oenb[5] la_oenb[60] la_oenb[61]
+ la_oenb[62] la_oenb[63] la_oenb[64] la_oenb[65] la_oenb[66] la_oenb[67] la_oenb[68]
+ la_oenb[69] la_oenb[6] la_oenb[70] la_oenb[71] la_oenb[72] la_oenb[73] la_oenb[74]
+ la_oenb[75] la_oenb[76] la_oenb[77] la_oenb[78] la_oenb[79] la_oenb[7] la_oenb[80]
+ la_oenb[81] la_oenb[82] la_oenb[83] la_oenb[84] la_oenb[85] la_oenb[86] la_oenb[87]
+ la_oenb[88] la_oenb[89] la_oenb[8] la_oenb[90] la_oenb[91] la_oenb[92] la_oenb[93]
+ la_oenb[94] la_oenb[95] la_oenb[96] la_oenb[97] la_oenb[98] la_oenb[99] la_oenb[9]
+ load_data load_status[0] load_status[1] load_status[2] master_ena_proc next_key
+ slv_done trigLoad vccd1 vssd1 wb_clk_i wb_rst_i
.ends

.subckt user_project_wrapper analog_io[0] analog_io[10] analog_io[11] analog_io[12]
+ analog_io[13] analog_io[14] analog_io[15] analog_io[16] analog_io[17] analog_io[18]
+ analog_io[19] analog_io[1] analog_io[20] analog_io[21] analog_io[22] analog_io[23]
+ analog_io[24] analog_io[25] analog_io[26] analog_io[27] analog_io[28] analog_io[2]
+ analog_io[3] analog_io[4] analog_io[5] analog_io[6] analog_io[7] analog_io[8] analog_io[9]
+ io_in[0] io_in[10] io_in[11] io_in[12] io_in[13] io_in[14] io_in[15] io_in[16] io_in[17]
+ io_in[18] io_in[19] io_in[1] io_in[20] io_in[21] io_in[22] io_in[23] io_in[24] io_in[25]
+ io_in[26] io_in[27] io_in[28] io_in[29] io_in[2] io_in[30] io_in[31] io_in[32] io_in[33]
+ io_in[34] io_in[35] io_in[36] io_in[37] io_in[3] io_in[4] io_in[5] io_in[6] io_in[7]
+ io_in[8] io_in[9] io_oeb[0] io_oeb[10] io_oeb[11] io_oeb[12] io_oeb[13] io_oeb[14]
+ io_oeb[15] io_oeb[16] io_oeb[17] io_oeb[18] io_oeb[19] io_oeb[1] io_oeb[20] io_oeb[21]
+ io_oeb[22] io_oeb[23] io_oeb[24] io_oeb[25] io_oeb[26] io_oeb[27] io_oeb[28] io_oeb[29]
+ io_oeb[2] io_oeb[30] io_oeb[31] io_oeb[32] io_oeb[33] io_oeb[34] io_oeb[35] io_oeb[36]
+ io_oeb[37] io_oeb[3] io_oeb[4] io_oeb[5] io_oeb[6] io_oeb[7] io_oeb[8] io_oeb[9]
+ io_out[0] io_out[10] io_out[11] io_out[12] io_out[13] io_out[14] io_out[15] io_out[16]
+ io_out[17] io_out[18] io_out[19] io_out[1] io_out[20] io_out[21] io_out[22] io_out[23]
+ io_out[24] io_out[25] io_out[26] io_out[27] io_out[28] io_out[29] io_out[2] io_out[30]
+ io_out[31] io_out[32] io_out[33] io_out[34] io_out[35] io_out[36] io_out[37] io_out[3]
+ io_out[4] io_out[5] io_out[6] io_out[7] io_out[8] io_out[9] la_data_in[0] la_data_in[100]
+ la_data_in[101] la_data_in[102] la_data_in[103] la_data_in[104] la_data_in[105]
+ la_data_in[106] la_data_in[107] la_data_in[108] la_data_in[109] la_data_in[10] la_data_in[110]
+ la_data_in[111] la_data_in[112] la_data_in[113] la_data_in[114] la_data_in[115]
+ la_data_in[116] la_data_in[117] la_data_in[118] la_data_in[119] la_data_in[11] la_data_in[120]
+ la_data_in[121] la_data_in[122] la_data_in[123] la_data_in[124] la_data_in[125]
+ la_data_in[126] la_data_in[127] la_data_in[12] la_data_in[13] la_data_in[14] la_data_in[15]
+ la_data_in[16] la_data_in[17] la_data_in[18] la_data_in[19] la_data_in[1] la_data_in[20]
+ la_data_in[21] la_data_in[22] la_data_in[23] la_data_in[24] la_data_in[25] la_data_in[26]
+ la_data_in[27] la_data_in[28] la_data_in[29] la_data_in[2] la_data_in[30] la_data_in[31]
+ la_data_in[32] la_data_in[33] la_data_in[34] la_data_in[35] la_data_in[36] la_data_in[37]
+ la_data_in[38] la_data_in[39] la_data_in[3] la_data_in[40] la_data_in[41] la_data_in[42]
+ la_data_in[43] la_data_in[44] la_data_in[45] la_data_in[46] la_data_in[47] la_data_in[48]
+ la_data_in[49] la_data_in[4] la_data_in[50] la_data_in[51] la_data_in[52] la_data_in[53]
+ la_data_in[54] la_data_in[55] la_data_in[56] la_data_in[57] la_data_in[58] la_data_in[59]
+ la_data_in[5] la_data_in[60] la_data_in[61] la_data_in[62] la_data_in[63] la_data_in[64]
+ la_data_in[65] la_data_in[66] la_data_in[67] la_data_in[68] la_data_in[69] la_data_in[6]
+ la_data_in[70] la_data_in[71] la_data_in[72] la_data_in[73] la_data_in[74] la_data_in[75]
+ la_data_in[76] la_data_in[77] la_data_in[78] la_data_in[79] la_data_in[7] la_data_in[80]
+ la_data_in[81] la_data_in[82] la_data_in[83] la_data_in[84] la_data_in[85] la_data_in[86]
+ la_data_in[87] la_data_in[88] la_data_in[89] la_data_in[8] la_data_in[90] la_data_in[91]
+ la_data_in[92] la_data_in[93] la_data_in[94] la_data_in[95] la_data_in[96] la_data_in[97]
+ la_data_in[98] la_data_in[99] la_data_in[9] la_data_out[0] la_data_out[100] la_data_out[101]
+ la_data_out[102] la_data_out[103] la_data_out[104] la_data_out[105] la_data_out[106]
+ la_data_out[107] la_data_out[108] la_data_out[109] la_data_out[10] la_data_out[110]
+ la_data_out[111] la_data_out[112] la_data_out[113] la_data_out[114] la_data_out[115]
+ la_data_out[116] la_data_out[117] la_data_out[118] la_data_out[119] la_data_out[11]
+ la_data_out[120] la_data_out[121] la_data_out[122] la_data_out[123] la_data_out[124]
+ la_data_out[125] la_data_out[126] la_data_out[127] la_data_out[12] la_data_out[13]
+ la_data_out[14] la_data_out[15] la_data_out[16] la_data_out[17] la_data_out[18]
+ la_data_out[19] la_data_out[1] la_data_out[20] la_data_out[21] la_data_out[22] la_data_out[23]
+ la_data_out[24] la_data_out[25] la_data_out[26] la_data_out[27] la_data_out[28]
+ la_data_out[29] la_data_out[2] la_data_out[30] la_data_out[31] la_data_out[32] la_data_out[33]
+ la_data_out[34] la_data_out[35] la_data_out[36] la_data_out[37] la_data_out[38]
+ la_data_out[39] la_data_out[3] la_data_out[40] la_data_out[41] la_data_out[42] la_data_out[43]
+ la_data_out[44] la_data_out[45] la_data_out[46] la_data_out[47] la_data_out[48]
+ la_data_out[49] la_data_out[4] la_data_out[50] la_data_out[51] la_data_out[52] la_data_out[53]
+ la_data_out[54] la_data_out[55] la_data_out[56] la_data_out[57] la_data_out[58]
+ la_data_out[59] la_data_out[5] la_data_out[60] la_data_out[61] la_data_out[62] la_data_out[63]
+ la_data_out[64] la_data_out[65] la_data_out[66] la_data_out[67] la_data_out[68]
+ la_data_out[69] la_data_out[6] la_data_out[70] la_data_out[71] la_data_out[72] la_data_out[73]
+ la_data_out[74] la_data_out[75] la_data_out[76] la_data_out[77] la_data_out[78]
+ la_data_out[79] la_data_out[7] la_data_out[80] la_data_out[81] la_data_out[82] la_data_out[83]
+ la_data_out[84] la_data_out[85] la_data_out[86] la_data_out[87] la_data_out[88]
+ la_data_out[89] la_data_out[8] la_data_out[90] la_data_out[91] la_data_out[92] la_data_out[93]
+ la_data_out[94] la_data_out[95] la_data_out[96] la_data_out[97] la_data_out[98]
+ la_data_out[99] la_data_out[9] la_oenb[0] la_oenb[100] la_oenb[101] la_oenb[102]
+ la_oenb[103] la_oenb[104] la_oenb[105] la_oenb[106] la_oenb[107] la_oenb[108] la_oenb[109]
+ la_oenb[10] la_oenb[110] la_oenb[111] la_oenb[112] la_oenb[113] la_oenb[114] la_oenb[115]
+ la_oenb[116] la_oenb[117] la_oenb[118] la_oenb[119] la_oenb[11] la_oenb[120] la_oenb[121]
+ la_oenb[122] la_oenb[123] la_oenb[124] la_oenb[125] la_oenb[126] la_oenb[127] la_oenb[12]
+ la_oenb[13] la_oenb[14] la_oenb[15] la_oenb[16] la_oenb[17] la_oenb[18] la_oenb[19]
+ la_oenb[1] la_oenb[20] la_oenb[21] la_oenb[22] la_oenb[23] la_oenb[24] la_oenb[25]
+ la_oenb[26] la_oenb[27] la_oenb[28] la_oenb[29] la_oenb[2] la_oenb[30] la_oenb[31]
+ la_oenb[32] la_oenb[33] la_oenb[34] la_oenb[35] la_oenb[36] la_oenb[37] la_oenb[38]
+ la_oenb[39] la_oenb[3] la_oenb[40] la_oenb[41] la_oenb[42] la_oenb[43] la_oenb[44]
+ la_oenb[45] la_oenb[46] la_oenb[47] la_oenb[48] la_oenb[49] la_oenb[4] la_oenb[50]
+ la_oenb[51] la_oenb[52] la_oenb[53] la_oenb[54] la_oenb[55] la_oenb[56] la_oenb[57]
+ la_oenb[58] la_oenb[59] la_oenb[5] la_oenb[60] la_oenb[61] la_oenb[62] la_oenb[63]
+ la_oenb[64] la_oenb[65] la_oenb[66] la_oenb[67] la_oenb[68] la_oenb[69] la_oenb[6]
+ la_oenb[70] la_oenb[71] la_oenb[72] la_oenb[73] la_oenb[74] la_oenb[75] la_oenb[76]
+ la_oenb[77] la_oenb[78] la_oenb[79] la_oenb[7] la_oenb[80] la_oenb[81] la_oenb[82]
+ la_oenb[83] la_oenb[84] la_oenb[85] la_oenb[86] la_oenb[87] la_oenb[88] la_oenb[89]
+ la_oenb[8] la_oenb[90] la_oenb[91] la_oenb[92] la_oenb[93] la_oenb[94] la_oenb[95]
+ la_oenb[96] la_oenb[97] la_oenb[98] la_oenb[99] la_oenb[9] user_clock2 user_irq[0]
+ user_irq[1] user_irq[2] vccd1 vccd2 vdda1 vdda2 vssa1 vssa2 vssd1 vssd2 wb_clk_i
+ wb_rst_i wbs_ack_o wbs_adr_i[0] wbs_adr_i[10] wbs_adr_i[11] wbs_adr_i[12] wbs_adr_i[13]
+ wbs_adr_i[14] wbs_adr_i[15] wbs_adr_i[16] wbs_adr_i[17] wbs_adr_i[18] wbs_adr_i[19]
+ wbs_adr_i[1] wbs_adr_i[20] wbs_adr_i[21] wbs_adr_i[22] wbs_adr_i[23] wbs_adr_i[24]
+ wbs_adr_i[25] wbs_adr_i[26] wbs_adr_i[27] wbs_adr_i[28] wbs_adr_i[29] wbs_adr_i[2]
+ wbs_adr_i[30] wbs_adr_i[31] wbs_adr_i[3] wbs_adr_i[4] wbs_adr_i[5] wbs_adr_i[6]
+ wbs_adr_i[7] wbs_adr_i[8] wbs_adr_i[9] wbs_cyc_i wbs_dat_i[0] wbs_dat_i[10] wbs_dat_i[11]
+ wbs_dat_i[12] wbs_dat_i[13] wbs_dat_i[14] wbs_dat_i[15] wbs_dat_i[16] wbs_dat_i[17]
+ wbs_dat_i[18] wbs_dat_i[19] wbs_dat_i[1] wbs_dat_i[20] wbs_dat_i[21] wbs_dat_i[22]
+ wbs_dat_i[23] wbs_dat_i[24] wbs_dat_i[25] wbs_dat_i[26] wbs_dat_i[27] wbs_dat_i[28]
+ wbs_dat_i[29] wbs_dat_i[2] wbs_dat_i[30] wbs_dat_i[31] wbs_dat_i[3] wbs_dat_i[4]
+ wbs_dat_i[5] wbs_dat_i[6] wbs_dat_i[7] wbs_dat_i[8] wbs_dat_i[9] wbs_dat_o[0] wbs_dat_o[10]
+ wbs_dat_o[11] wbs_dat_o[12] wbs_dat_o[13] wbs_dat_o[14] wbs_dat_o[15] wbs_dat_o[16]
+ wbs_dat_o[17] wbs_dat_o[18] wbs_dat_o[19] wbs_dat_o[1] wbs_dat_o[20] wbs_dat_o[21]
+ wbs_dat_o[22] wbs_dat_o[23] wbs_dat_o[24] wbs_dat_o[25] wbs_dat_o[26] wbs_dat_o[27]
+ wbs_dat_o[28] wbs_dat_o[29] wbs_dat_o[2] wbs_dat_o[30] wbs_dat_o[31] wbs_dat_o[3]
+ wbs_dat_o[4] wbs_dat_o[5] wbs_dat_o[6] wbs_dat_o[7] wbs_dat_o[8] wbs_dat_o[9] wbs_sel_i[0]
+ wbs_sel_i[1] wbs_sel_i[2] wbs_sel_i[3] wbs_stb_i wbs_we_i
Xbec_core bec_core/becStatus[0] bec_core/becStatus[1] bec_core/becStatus[2] bec_core/becStatus[3]
+ wb_clk_i bec_core/data_in[0] bec_core/data_in[100] bec_core/data_in[101] bec_core/data_in[102]
+ bec_core/data_in[103] bec_core/data_in[104] bec_core/data_in[105] bec_core/data_in[106]
+ bec_core/data_in[107] bec_core/data_in[108] bec_core/data_in[109] bec_core/data_in[10]
+ bec_core/data_in[110] bec_core/data_in[111] bec_core/data_in[112] bec_core/data_in[113]
+ bec_core/data_in[114] bec_core/data_in[115] bec_core/data_in[116] bec_core/data_in[117]
+ bec_core/data_in[118] bec_core/data_in[119] bec_core/data_in[11] bec_core/data_in[120]
+ bec_core/data_in[121] bec_core/data_in[122] bec_core/data_in[123] bec_core/data_in[124]
+ bec_core/data_in[125] bec_core/data_in[126] bec_core/data_in[127] bec_core/data_in[128]
+ bec_core/data_in[129] bec_core/data_in[12] bec_core/data_in[130] bec_core/data_in[131]
+ bec_core/data_in[132] bec_core/data_in[133] bec_core/data_in[134] bec_core/data_in[135]
+ bec_core/data_in[136] bec_core/data_in[137] bec_core/data_in[138] bec_core/data_in[139]
+ bec_core/data_in[13] bec_core/data_in[140] bec_core/data_in[141] bec_core/data_in[142]
+ bec_core/data_in[143] bec_core/data_in[144] bec_core/data_in[145] bec_core/data_in[146]
+ bec_core/data_in[147] bec_core/data_in[148] bec_core/data_in[149] bec_core/data_in[14]
+ bec_core/data_in[150] bec_core/data_in[151] bec_core/data_in[152] bec_core/data_in[153]
+ bec_core/data_in[154] bec_core/data_in[155] bec_core/data_in[156] bec_core/data_in[157]
+ bec_core/data_in[158] bec_core/data_in[159] bec_core/data_in[15] bec_core/data_in[160]
+ bec_core/data_in[161] bec_core/data_in[162] bec_core/data_in[16] bec_core/data_in[17]
+ bec_core/data_in[18] bec_core/data_in[19] bec_core/data_in[1] bec_core/data_in[20]
+ bec_core/data_in[21] bec_core/data_in[22] bec_core/data_in[23] bec_core/data_in[24]
+ bec_core/data_in[25] bec_core/data_in[26] bec_core/data_in[27] bec_core/data_in[28]
+ bec_core/data_in[29] bec_core/data_in[2] bec_core/data_in[30] bec_core/data_in[31]
+ bec_core/data_in[32] bec_core/data_in[33] bec_core/data_in[34] bec_core/data_in[35]
+ bec_core/data_in[36] bec_core/data_in[37] bec_core/data_in[38] bec_core/data_in[39]
+ bec_core/data_in[3] bec_core/data_in[40] bec_core/data_in[41] bec_core/data_in[42]
+ bec_core/data_in[43] bec_core/data_in[44] bec_core/data_in[45] bec_core/data_in[46]
+ bec_core/data_in[47] bec_core/data_in[48] bec_core/data_in[49] bec_core/data_in[4]
+ bec_core/data_in[50] bec_core/data_in[51] bec_core/data_in[52] bec_core/data_in[53]
+ bec_core/data_in[54] bec_core/data_in[55] bec_core/data_in[56] bec_core/data_in[57]
+ bec_core/data_in[58] bec_core/data_in[59] bec_core/data_in[5] bec_core/data_in[60]
+ bec_core/data_in[61] bec_core/data_in[62] bec_core/data_in[63] bec_core/data_in[64]
+ bec_core/data_in[65] bec_core/data_in[66] bec_core/data_in[67] bec_core/data_in[68]
+ bec_core/data_in[69] bec_core/data_in[6] bec_core/data_in[70] bec_core/data_in[71]
+ bec_core/data_in[72] bec_core/data_in[73] bec_core/data_in[74] bec_core/data_in[75]
+ bec_core/data_in[76] bec_core/data_in[77] bec_core/data_in[78] bec_core/data_in[79]
+ bec_core/data_in[7] bec_core/data_in[80] bec_core/data_in[81] bec_core/data_in[82]
+ bec_core/data_in[83] bec_core/data_in[84] bec_core/data_in[85] bec_core/data_in[86]
+ bec_core/data_in[87] bec_core/data_in[88] bec_core/data_in[89] bec_core/data_in[8]
+ bec_core/data_in[90] bec_core/data_in[91] bec_core/data_in[92] bec_core/data_in[93]
+ bec_core/data_in[94] bec_core/data_in[95] bec_core/data_in[96] bec_core/data_in[97]
+ bec_core/data_in[98] bec_core/data_in[99] bec_core/data_in[9] bec_core/data_out[0]
+ bec_core/data_out[100] bec_core/data_out[101] bec_core/data_out[102] bec_core/data_out[103]
+ bec_core/data_out[104] bec_core/data_out[105] bec_core/data_out[106] bec_core/data_out[107]
+ bec_core/data_out[108] bec_core/data_out[109] bec_core/data_out[10] bec_core/data_out[110]
+ bec_core/data_out[111] bec_core/data_out[112] bec_core/data_out[113] bec_core/data_out[114]
+ bec_core/data_out[115] bec_core/data_out[116] bec_core/data_out[117] bec_core/data_out[118]
+ bec_core/data_out[119] bec_core/data_out[11] bec_core/data_out[120] bec_core/data_out[121]
+ bec_core/data_out[122] bec_core/data_out[123] bec_core/data_out[124] bec_core/data_out[125]
+ bec_core/data_out[126] bec_core/data_out[127] bec_core/data_out[128] bec_core/data_out[129]
+ bec_core/data_out[12] bec_core/data_out[130] bec_core/data_out[131] bec_core/data_out[132]
+ bec_core/data_out[133] bec_core/data_out[134] bec_core/data_out[135] bec_core/data_out[136]
+ bec_core/data_out[137] bec_core/data_out[138] bec_core/data_out[139] bec_core/data_out[13]
+ bec_core/data_out[140] bec_core/data_out[141] bec_core/data_out[142] bec_core/data_out[143]
+ bec_core/data_out[144] bec_core/data_out[145] bec_core/data_out[146] bec_core/data_out[147]
+ bec_core/data_out[148] bec_core/data_out[149] bec_core/data_out[14] bec_core/data_out[150]
+ bec_core/data_out[151] bec_core/data_out[152] bec_core/data_out[153] bec_core/data_out[154]
+ bec_core/data_out[155] bec_core/data_out[156] bec_core/data_out[157] bec_core/data_out[158]
+ bec_core/data_out[159] bec_core/data_out[15] bec_core/data_out[160] bec_core/data_out[161]
+ bec_core/data_out[162] bec_core/data_out[16] bec_core/data_out[17] bec_core/data_out[18]
+ bec_core/data_out[19] bec_core/data_out[1] bec_core/data_out[20] bec_core/data_out[21]
+ bec_core/data_out[22] bec_core/data_out[23] bec_core/data_out[24] bec_core/data_out[25]
+ bec_core/data_out[26] bec_core/data_out[27] bec_core/data_out[28] bec_core/data_out[29]
+ bec_core/data_out[2] bec_core/data_out[30] bec_core/data_out[31] bec_core/data_out[32]
+ bec_core/data_out[33] bec_core/data_out[34] bec_core/data_out[35] bec_core/data_out[36]
+ bec_core/data_out[37] bec_core/data_out[38] bec_core/data_out[39] bec_core/data_out[3]
+ bec_core/data_out[40] bec_core/data_out[41] bec_core/data_out[42] bec_core/data_out[43]
+ bec_core/data_out[44] bec_core/data_out[45] bec_core/data_out[46] bec_core/data_out[47]
+ bec_core/data_out[48] bec_core/data_out[49] bec_core/data_out[4] bec_core/data_out[50]
+ bec_core/data_out[51] bec_core/data_out[52] bec_core/data_out[53] bec_core/data_out[54]
+ bec_core/data_out[55] bec_core/data_out[56] bec_core/data_out[57] bec_core/data_out[58]
+ bec_core/data_out[59] bec_core/data_out[5] bec_core/data_out[60] bec_core/data_out[61]
+ bec_core/data_out[62] bec_core/data_out[63] bec_core/data_out[64] bec_core/data_out[65]
+ bec_core/data_out[66] bec_core/data_out[67] bec_core/data_out[68] bec_core/data_out[69]
+ bec_core/data_out[6] bec_core/data_out[70] bec_core/data_out[71] bec_core/data_out[72]
+ bec_core/data_out[73] bec_core/data_out[74] bec_core/data_out[75] bec_core/data_out[76]
+ bec_core/data_out[77] bec_core/data_out[78] bec_core/data_out[79] bec_core/data_out[7]
+ bec_core/data_out[80] bec_core/data_out[81] bec_core/data_out[82] bec_core/data_out[83]
+ bec_core/data_out[84] bec_core/data_out[85] bec_core/data_out[86] bec_core/data_out[87]
+ bec_core/data_out[88] bec_core/data_out[89] bec_core/data_out[8] bec_core/data_out[90]
+ bec_core/data_out[91] bec_core/data_out[92] bec_core/data_out[93] bec_core/data_out[94]
+ bec_core/data_out[95] bec_core/data_out[96] bec_core/data_out[97] bec_core/data_out[98]
+ bec_core/data_out[99] bec_core/data_out[9] bec_core/done bec_core/enable bec_core/ki
+ bec_core/load_data bec_core/load_status[0] bec_core/load_status[1] bec_core/load_status[2]
+ bec_core/next_key wb_rst_i bec_core/trigLoad vccd2 vssd2 sm_bec_v3
Xcontrol_unit bec_core/becStatus[0] bec_core/becStatus[1] bec_core/becStatus[2] bec_core/becStatus[3]
+ bec_core/data_out[0] bec_core/data_out[100] bec_core/data_out[101] bec_core/data_out[102]
+ bec_core/data_out[103] bec_core/data_out[104] bec_core/data_out[105] bec_core/data_out[106]
+ bec_core/data_out[107] bec_core/data_out[108] bec_core/data_out[109] bec_core/data_out[10]
+ bec_core/data_out[110] bec_core/data_out[111] bec_core/data_out[112] bec_core/data_out[113]
+ bec_core/data_out[114] bec_core/data_out[115] bec_core/data_out[116] bec_core/data_out[117]
+ bec_core/data_out[118] bec_core/data_out[119] bec_core/data_out[11] bec_core/data_out[120]
+ bec_core/data_out[121] bec_core/data_out[122] bec_core/data_out[123] bec_core/data_out[124]
+ bec_core/data_out[125] bec_core/data_out[126] bec_core/data_out[127] bec_core/data_out[128]
+ bec_core/data_out[129] bec_core/data_out[12] bec_core/data_out[130] bec_core/data_out[131]
+ bec_core/data_out[132] bec_core/data_out[133] bec_core/data_out[134] bec_core/data_out[135]
+ bec_core/data_out[136] bec_core/data_out[137] bec_core/data_out[138] bec_core/data_out[139]
+ bec_core/data_out[13] bec_core/data_out[140] bec_core/data_out[141] bec_core/data_out[142]
+ bec_core/data_out[143] bec_core/data_out[144] bec_core/data_out[145] bec_core/data_out[146]
+ bec_core/data_out[147] bec_core/data_out[148] bec_core/data_out[149] bec_core/data_out[14]
+ bec_core/data_out[150] bec_core/data_out[151] bec_core/data_out[152] bec_core/data_out[153]
+ bec_core/data_out[154] bec_core/data_out[155] bec_core/data_out[156] bec_core/data_out[157]
+ bec_core/data_out[158] bec_core/data_out[159] bec_core/data_out[15] bec_core/data_out[160]
+ bec_core/data_out[161] bec_core/data_out[162] bec_core/data_out[16] bec_core/data_out[17]
+ bec_core/data_out[18] bec_core/data_out[19] bec_core/data_out[1] bec_core/data_out[20]
+ bec_core/data_out[21] bec_core/data_out[22] bec_core/data_out[23] bec_core/data_out[24]
+ bec_core/data_out[25] bec_core/data_out[26] bec_core/data_out[27] bec_core/data_out[28]
+ bec_core/data_out[29] bec_core/data_out[2] bec_core/data_out[30] bec_core/data_out[31]
+ bec_core/data_out[32] bec_core/data_out[33] bec_core/data_out[34] bec_core/data_out[35]
+ bec_core/data_out[36] bec_core/data_out[37] bec_core/data_out[38] bec_core/data_out[39]
+ bec_core/data_out[3] bec_core/data_out[40] bec_core/data_out[41] bec_core/data_out[42]
+ bec_core/data_out[43] bec_core/data_out[44] bec_core/data_out[45] bec_core/data_out[46]
+ bec_core/data_out[47] bec_core/data_out[48] bec_core/data_out[49] bec_core/data_out[4]
+ bec_core/data_out[50] bec_core/data_out[51] bec_core/data_out[52] bec_core/data_out[53]
+ bec_core/data_out[54] bec_core/data_out[55] bec_core/data_out[56] bec_core/data_out[57]
+ bec_core/data_out[58] bec_core/data_out[59] bec_core/data_out[5] bec_core/data_out[60]
+ bec_core/data_out[61] bec_core/data_out[62] bec_core/data_out[63] bec_core/data_out[64]
+ bec_core/data_out[65] bec_core/data_out[66] bec_core/data_out[67] bec_core/data_out[68]
+ bec_core/data_out[69] bec_core/data_out[6] bec_core/data_out[70] bec_core/data_out[71]
+ bec_core/data_out[72] bec_core/data_out[73] bec_core/data_out[74] bec_core/data_out[75]
+ bec_core/data_out[76] bec_core/data_out[77] bec_core/data_out[78] bec_core/data_out[79]
+ bec_core/data_out[7] bec_core/data_out[80] bec_core/data_out[81] bec_core/data_out[82]
+ bec_core/data_out[83] bec_core/data_out[84] bec_core/data_out[85] bec_core/data_out[86]
+ bec_core/data_out[87] bec_core/data_out[88] bec_core/data_out[89] bec_core/data_out[8]
+ bec_core/data_out[90] bec_core/data_out[91] bec_core/data_out[92] bec_core/data_out[93]
+ bec_core/data_out[94] bec_core/data_out[95] bec_core/data_out[96] bec_core/data_out[97]
+ bec_core/data_out[98] bec_core/data_out[99] bec_core/data_out[9] bec_core/data_in[0]
+ bec_core/data_in[100] bec_core/data_in[101] bec_core/data_in[102] bec_core/data_in[103]
+ bec_core/data_in[104] bec_core/data_in[105] bec_core/data_in[106] bec_core/data_in[107]
+ bec_core/data_in[108] bec_core/data_in[109] bec_core/data_in[10] bec_core/data_in[110]
+ bec_core/data_in[111] bec_core/data_in[112] bec_core/data_in[113] bec_core/data_in[114]
+ bec_core/data_in[115] bec_core/data_in[116] bec_core/data_in[117] bec_core/data_in[118]
+ bec_core/data_in[119] bec_core/data_in[11] bec_core/data_in[120] bec_core/data_in[121]
+ bec_core/data_in[122] bec_core/data_in[123] bec_core/data_in[124] bec_core/data_in[125]
+ bec_core/data_in[126] bec_core/data_in[127] bec_core/data_in[128] bec_core/data_in[129]
+ bec_core/data_in[12] bec_core/data_in[130] bec_core/data_in[131] bec_core/data_in[132]
+ bec_core/data_in[133] bec_core/data_in[134] bec_core/data_in[135] bec_core/data_in[136]
+ bec_core/data_in[137] bec_core/data_in[138] bec_core/data_in[139] bec_core/data_in[13]
+ bec_core/data_in[140] bec_core/data_in[141] bec_core/data_in[142] bec_core/data_in[143]
+ bec_core/data_in[144] bec_core/data_in[145] bec_core/data_in[146] bec_core/data_in[147]
+ bec_core/data_in[148] bec_core/data_in[149] bec_core/data_in[14] bec_core/data_in[150]
+ bec_core/data_in[151] bec_core/data_in[152] bec_core/data_in[153] bec_core/data_in[154]
+ bec_core/data_in[155] bec_core/data_in[156] bec_core/data_in[157] bec_core/data_in[158]
+ bec_core/data_in[159] bec_core/data_in[15] bec_core/data_in[160] bec_core/data_in[161]
+ bec_core/data_in[162] bec_core/data_in[16] bec_core/data_in[17] bec_core/data_in[18]
+ bec_core/data_in[19] bec_core/data_in[1] bec_core/data_in[20] bec_core/data_in[21]
+ bec_core/data_in[22] bec_core/data_in[23] bec_core/data_in[24] bec_core/data_in[25]
+ bec_core/data_in[26] bec_core/data_in[27] bec_core/data_in[28] bec_core/data_in[29]
+ bec_core/data_in[2] bec_core/data_in[30] bec_core/data_in[31] bec_core/data_in[32]
+ bec_core/data_in[33] bec_core/data_in[34] bec_core/data_in[35] bec_core/data_in[36]
+ bec_core/data_in[37] bec_core/data_in[38] bec_core/data_in[39] bec_core/data_in[3]
+ bec_core/data_in[40] bec_core/data_in[41] bec_core/data_in[42] bec_core/data_in[43]
+ bec_core/data_in[44] bec_core/data_in[45] bec_core/data_in[46] bec_core/data_in[47]
+ bec_core/data_in[48] bec_core/data_in[49] bec_core/data_in[4] bec_core/data_in[50]
+ bec_core/data_in[51] bec_core/data_in[52] bec_core/data_in[53] bec_core/data_in[54]
+ bec_core/data_in[55] bec_core/data_in[56] bec_core/data_in[57] bec_core/data_in[58]
+ bec_core/data_in[59] bec_core/data_in[5] bec_core/data_in[60] bec_core/data_in[61]
+ bec_core/data_in[62] bec_core/data_in[63] bec_core/data_in[64] bec_core/data_in[65]
+ bec_core/data_in[66] bec_core/data_in[67] bec_core/data_in[68] bec_core/data_in[69]
+ bec_core/data_in[6] bec_core/data_in[70] bec_core/data_in[71] bec_core/data_in[72]
+ bec_core/data_in[73] bec_core/data_in[74] bec_core/data_in[75] bec_core/data_in[76]
+ bec_core/data_in[77] bec_core/data_in[78] bec_core/data_in[79] bec_core/data_in[7]
+ bec_core/data_in[80] bec_core/data_in[81] bec_core/data_in[82] bec_core/data_in[83]
+ bec_core/data_in[84] bec_core/data_in[85] bec_core/data_in[86] bec_core/data_in[87]
+ bec_core/data_in[88] bec_core/data_in[89] bec_core/data_in[8] bec_core/data_in[90]
+ bec_core/data_in[91] bec_core/data_in[92] bec_core/data_in[93] bec_core/data_in[94]
+ bec_core/data_in[95] bec_core/data_in[96] bec_core/data_in[97] bec_core/data_in[98]
+ bec_core/data_in[99] bec_core/data_in[9] bec_core/ki la_data_in[0] la_data_in[100]
+ la_data_in[101] la_data_in[102] la_data_in[103] la_data_in[104] la_data_in[105]
+ la_data_in[106] la_data_in[107] la_data_in[108] la_data_in[109] la_data_in[10] la_data_in[110]
+ la_data_in[111] la_data_in[112] la_data_in[113] la_data_in[114] la_data_in[115]
+ la_data_in[116] la_data_in[117] la_data_in[118] la_data_in[119] la_data_in[11] la_data_in[120]
+ la_data_in[121] la_data_in[122] la_data_in[123] la_data_in[124] la_data_in[125]
+ la_data_in[126] la_data_in[127] la_data_in[12] la_data_in[13] la_data_in[14] la_data_in[15]
+ la_data_in[16] la_data_in[17] la_data_in[18] la_data_in[19] la_data_in[1] la_data_in[20]
+ la_data_in[21] la_data_in[22] la_data_in[23] la_data_in[24] la_data_in[25] la_data_in[26]
+ la_data_in[27] la_data_in[28] la_data_in[29] la_data_in[2] la_data_in[30] la_data_in[31]
+ la_data_in[32] la_data_in[33] la_data_in[34] la_data_in[35] la_data_in[36] la_data_in[37]
+ la_data_in[38] la_data_in[39] la_data_in[3] la_data_in[40] la_data_in[41] la_data_in[42]
+ la_data_in[43] la_data_in[44] la_data_in[45] la_data_in[46] la_data_in[47] la_data_in[48]
+ la_data_in[49] la_data_in[4] la_data_in[50] la_data_in[51] la_data_in[52] la_data_in[53]
+ la_data_in[54] la_data_in[55] la_data_in[56] la_data_in[57] la_data_in[58] la_data_in[59]
+ la_data_in[5] la_data_in[60] la_data_in[61] la_data_in[62] la_data_in[63] la_data_in[64]
+ la_data_in[65] la_data_in[66] la_data_in[67] la_data_in[68] la_data_in[69] la_data_in[6]
+ la_data_in[70] la_data_in[71] la_data_in[72] la_data_in[73] la_data_in[74] la_data_in[75]
+ la_data_in[76] la_data_in[77] la_data_in[78] la_data_in[79] la_data_in[7] la_data_in[80]
+ la_data_in[81] la_data_in[82] la_data_in[83] la_data_in[84] la_data_in[85] la_data_in[86]
+ la_data_in[87] la_data_in[88] la_data_in[89] la_data_in[8] la_data_in[90] la_data_in[91]
+ la_data_in[92] la_data_in[93] la_data_in[94] la_data_in[95] la_data_in[96] la_data_in[97]
+ la_data_in[98] la_data_in[99] la_data_in[9] la_data_out[0] la_data_out[100] la_data_out[101]
+ la_data_out[102] la_data_out[103] la_data_out[104] la_data_out[105] la_data_out[106]
+ la_data_out[107] la_data_out[108] la_data_out[109] la_data_out[10] la_data_out[110]
+ la_data_out[111] la_data_out[112] la_data_out[113] la_data_out[114] la_data_out[115]
+ la_data_out[116] la_data_out[117] la_data_out[118] la_data_out[119] la_data_out[11]
+ la_data_out[120] la_data_out[121] la_data_out[122] la_data_out[123] la_data_out[124]
+ la_data_out[125] la_data_out[126] la_data_out[127] la_data_out[12] la_data_out[13]
+ la_data_out[14] la_data_out[15] la_data_out[16] la_data_out[17] la_data_out[18]
+ la_data_out[19] la_data_out[1] la_data_out[20] la_data_out[21] la_data_out[22] la_data_out[23]
+ la_data_out[24] la_data_out[25] la_data_out[26] la_data_out[27] la_data_out[28]
+ la_data_out[29] la_data_out[2] la_data_out[30] la_data_out[31] la_data_out[32] la_data_out[33]
+ la_data_out[34] la_data_out[35] la_data_out[36] la_data_out[37] la_data_out[38]
+ la_data_out[39] la_data_out[3] la_data_out[40] la_data_out[41] la_data_out[42] la_data_out[43]
+ la_data_out[44] la_data_out[45] la_data_out[46] la_data_out[47] la_data_out[48]
+ la_data_out[49] la_data_out[4] la_data_out[50] la_data_out[51] la_data_out[52] la_data_out[53]
+ la_data_out[54] la_data_out[55] la_data_out[56] la_data_out[57] la_data_out[58]
+ la_data_out[59] la_data_out[5] la_data_out[60] la_data_out[61] la_data_out[62] la_data_out[63]
+ la_data_out[64] la_data_out[65] la_data_out[66] la_data_out[67] la_data_out[68]
+ la_data_out[69] la_data_out[6] la_data_out[70] la_data_out[71] la_data_out[72] la_data_out[73]
+ la_data_out[74] la_data_out[75] la_data_out[76] la_data_out[77] la_data_out[78]
+ la_data_out[79] la_data_out[7] la_data_out[80] la_data_out[81] la_data_out[82] la_data_out[83]
+ la_data_out[84] la_data_out[85] la_data_out[86] la_data_out[87] la_data_out[88]
+ la_data_out[89] la_data_out[8] la_data_out[90] la_data_out[91] la_data_out[92] la_data_out[93]
+ la_data_out[94] la_data_out[95] la_data_out[96] la_data_out[97] la_data_out[98]
+ la_data_out[99] la_data_out[9] la_oenb[0] la_oenb[100] la_oenb[101] la_oenb[102]
+ la_oenb[103] la_oenb[104] la_oenb[105] la_oenb[106] la_oenb[107] la_oenb[108] la_oenb[109]
+ la_oenb[10] la_oenb[110] la_oenb[111] la_oenb[112] la_oenb[113] la_oenb[114] la_oenb[115]
+ la_oenb[116] la_oenb[117] la_oenb[118] la_oenb[119] la_oenb[11] la_oenb[120] la_oenb[121]
+ la_oenb[122] la_oenb[123] la_oenb[124] la_oenb[125] la_oenb[126] la_oenb[127] la_oenb[12]
+ la_oenb[13] la_oenb[14] la_oenb[15] la_oenb[16] la_oenb[17] la_oenb[18] la_oenb[19]
+ la_oenb[1] la_oenb[20] la_oenb[21] la_oenb[22] la_oenb[23] la_oenb[24] la_oenb[25]
+ la_oenb[26] la_oenb[27] la_oenb[28] la_oenb[29] la_oenb[2] la_oenb[30] la_oenb[31]
+ la_oenb[32] la_oenb[33] la_oenb[34] la_oenb[35] la_oenb[36] la_oenb[37] la_oenb[38]
+ la_oenb[39] la_oenb[3] la_oenb[40] la_oenb[41] la_oenb[42] la_oenb[43] la_oenb[44]
+ la_oenb[45] la_oenb[46] la_oenb[47] la_oenb[48] la_oenb[49] la_oenb[4] la_oenb[50]
+ la_oenb[51] la_oenb[52] la_oenb[53] la_oenb[54] la_oenb[55] la_oenb[56] la_oenb[57]
+ la_oenb[58] la_oenb[59] la_oenb[5] la_oenb[60] la_oenb[61] la_oenb[62] la_oenb[63]
+ la_oenb[64] la_oenb[65] la_oenb[66] la_oenb[67] la_oenb[68] la_oenb[69] la_oenb[6]
+ la_oenb[70] la_oenb[71] la_oenb[72] la_oenb[73] la_oenb[74] la_oenb[75] la_oenb[76]
+ la_oenb[77] la_oenb[78] la_oenb[79] la_oenb[7] la_oenb[80] la_oenb[81] la_oenb[82]
+ la_oenb[83] la_oenb[84] la_oenb[85] la_oenb[86] la_oenb[87] la_oenb[88] la_oenb[89]
+ la_oenb[8] la_oenb[90] la_oenb[91] la_oenb[92] la_oenb[93] la_oenb[94] la_oenb[95]
+ la_oenb[96] la_oenb[97] la_oenb[98] la_oenb[99] la_oenb[9] bec_core/load_data bec_core/load_status[0]
+ bec_core/load_status[1] bec_core/load_status[2] bec_core/enable bec_core/next_key
+ bec_core/done bec_core/trigLoad vccd1 vssd1 wb_clk_i wb_rst_i controller
.ends

