// This is the unpowered netlist.
module user_project_wrapper (user_clock2,
    wb_clk_i,
    wb_rst_i,
    wbs_ack_o,
    wbs_cyc_i,
    wbs_stb_i,
    wbs_we_i,
    analog_io,
    io_in,
    io_oeb,
    io_out,
    la_data_in,
    la_data_out,
    la_oenb,
    user_irq,
    wbs_adr_i,
    wbs_dat_i,
    wbs_dat_o,
    wbs_sel_i);
 input user_clock2;
 input wb_clk_i;
 input wb_rst_i;
 output wbs_ack_o;
 input wbs_cyc_i;
 input wbs_stb_i;
 input wbs_we_i;
 inout [28:0] analog_io;
 input [37:0] io_in;
 output [37:0] io_oeb;
 output [37:0] io_out;
 input [127:0] la_data_in;
 output [127:0] la_data_out;
 input [127:0] la_oenb;
 output [2:0] user_irq;
 input [31:0] wbs_adr_i;
 input [31:0] wbs_dat_i;
 output [31:0] wbs_dat_o;
 input [3:0] wbs_sel_i;

 wire \configBus[0] ;
 wire \configBus[100] ;
 wire \configBus[101] ;
 wire \configBus[102] ;
 wire \configBus[103] ;
 wire \configBus[104] ;
 wire \configBus[105] ;
 wire \configBus[106] ;
 wire \configBus[107] ;
 wire \configBus[108] ;
 wire \configBus[109] ;
 wire \configBus[10] ;
 wire \configBus[110] ;
 wire \configBus[111] ;
 wire \configBus[112] ;
 wire \configBus[113] ;
 wire \configBus[114] ;
 wire \configBus[115] ;
 wire \configBus[116] ;
 wire \configBus[117] ;
 wire \configBus[118] ;
 wire \configBus[119] ;
 wire \configBus[11] ;
 wire \configBus[120] ;
 wire \configBus[121] ;
 wire \configBus[122] ;
 wire \configBus[123] ;
 wire \configBus[124] ;
 wire \configBus[125] ;
 wire \configBus[126] ;
 wire \configBus[127] ;
 wire \configBus[128] ;
 wire \configBus[129] ;
 wire \configBus[12] ;
 wire \configBus[130] ;
 wire \configBus[131] ;
 wire \configBus[132] ;
 wire \configBus[133] ;
 wire \configBus[134] ;
 wire \configBus[135] ;
 wire \configBus[136] ;
 wire \configBus[137] ;
 wire \configBus[138] ;
 wire \configBus[139] ;
 wire \configBus[13] ;
 wire \configBus[140] ;
 wire \configBus[141] ;
 wire \configBus[142] ;
 wire \configBus[143] ;
 wire \configBus[144] ;
 wire \configBus[145] ;
 wire \configBus[146] ;
 wire \configBus[147] ;
 wire \configBus[148] ;
 wire \configBus[149] ;
 wire \configBus[14] ;
 wire \configBus[150] ;
 wire \configBus[151] ;
 wire \configBus[152] ;
 wire \configBus[153] ;
 wire \configBus[154] ;
 wire \configBus[155] ;
 wire \configBus[156] ;
 wire \configBus[157] ;
 wire \configBus[158] ;
 wire \configBus[159] ;
 wire \configBus[15] ;
 wire \configBus[160] ;
 wire \configBus[161] ;
 wire \configBus[162] ;
 wire \configBus[16] ;
 wire \configBus[17] ;
 wire \configBus[18] ;
 wire \configBus[19] ;
 wire \configBus[1] ;
 wire \configBus[20] ;
 wire \configBus[21] ;
 wire \configBus[22] ;
 wire \configBus[23] ;
 wire \configBus[24] ;
 wire \configBus[25] ;
 wire \configBus[26] ;
 wire \configBus[27] ;
 wire \configBus[28] ;
 wire \configBus[29] ;
 wire \configBus[2] ;
 wire \configBus[30] ;
 wire \configBus[31] ;
 wire \configBus[32] ;
 wire \configBus[33] ;
 wire \configBus[34] ;
 wire \configBus[35] ;
 wire \configBus[36] ;
 wire \configBus[37] ;
 wire \configBus[38] ;
 wire \configBus[39] ;
 wire \configBus[3] ;
 wire \configBus[40] ;
 wire \configBus[41] ;
 wire \configBus[42] ;
 wire \configBus[43] ;
 wire \configBus[44] ;
 wire \configBus[45] ;
 wire \configBus[46] ;
 wire \configBus[47] ;
 wire \configBus[48] ;
 wire \configBus[49] ;
 wire \configBus[4] ;
 wire \configBus[50] ;
 wire \configBus[51] ;
 wire \configBus[52] ;
 wire \configBus[53] ;
 wire \configBus[54] ;
 wire \configBus[55] ;
 wire \configBus[56] ;
 wire \configBus[57] ;
 wire \configBus[58] ;
 wire \configBus[59] ;
 wire \configBus[5] ;
 wire \configBus[60] ;
 wire \configBus[61] ;
 wire \configBus[62] ;
 wire \configBus[63] ;
 wire \configBus[64] ;
 wire \configBus[65] ;
 wire \configBus[66] ;
 wire \configBus[67] ;
 wire \configBus[68] ;
 wire \configBus[69] ;
 wire \configBus[6] ;
 wire \configBus[70] ;
 wire \configBus[71] ;
 wire \configBus[72] ;
 wire \configBus[73] ;
 wire \configBus[74] ;
 wire \configBus[75] ;
 wire \configBus[76] ;
 wire \configBus[77] ;
 wire \configBus[78] ;
 wire \configBus[79] ;
 wire \configBus[7] ;
 wire \configBus[80] ;
 wire \configBus[81] ;
 wire \configBus[82] ;
 wire \configBus[83] ;
 wire \configBus[84] ;
 wire \configBus[85] ;
 wire \configBus[86] ;
 wire \configBus[87] ;
 wire \configBus[88] ;
 wire \configBus[89] ;
 wire \configBus[8] ;
 wire \configBus[90] ;
 wire \configBus[91] ;
 wire \configBus[92] ;
 wire \configBus[93] ;
 wire \configBus[94] ;
 wire \configBus[95] ;
 wire \configBus[96] ;
 wire \configBus[97] ;
 wire \configBus[98] ;
 wire \configBus[99] ;
 wire \configBus[9] ;
 wire \dataBus[0] ;
 wire \dataBus[100] ;
 wire \dataBus[101] ;
 wire \dataBus[102] ;
 wire \dataBus[103] ;
 wire \dataBus[104] ;
 wire \dataBus[105] ;
 wire \dataBus[106] ;
 wire \dataBus[107] ;
 wire \dataBus[108] ;
 wire \dataBus[109] ;
 wire \dataBus[10] ;
 wire \dataBus[110] ;
 wire \dataBus[111] ;
 wire \dataBus[112] ;
 wire \dataBus[113] ;
 wire \dataBus[114] ;
 wire \dataBus[115] ;
 wire \dataBus[116] ;
 wire \dataBus[117] ;
 wire \dataBus[118] ;
 wire \dataBus[119] ;
 wire \dataBus[11] ;
 wire \dataBus[120] ;
 wire \dataBus[121] ;
 wire \dataBus[122] ;
 wire \dataBus[123] ;
 wire \dataBus[124] ;
 wire \dataBus[125] ;
 wire \dataBus[126] ;
 wire \dataBus[127] ;
 wire \dataBus[128] ;
 wire \dataBus[129] ;
 wire \dataBus[12] ;
 wire \dataBus[130] ;
 wire \dataBus[131] ;
 wire \dataBus[132] ;
 wire \dataBus[133] ;
 wire \dataBus[134] ;
 wire \dataBus[135] ;
 wire \dataBus[136] ;
 wire \dataBus[137] ;
 wire \dataBus[138] ;
 wire \dataBus[139] ;
 wire \dataBus[13] ;
 wire \dataBus[140] ;
 wire \dataBus[141] ;
 wire \dataBus[142] ;
 wire \dataBus[143] ;
 wire \dataBus[144] ;
 wire \dataBus[145] ;
 wire \dataBus[146] ;
 wire \dataBus[147] ;
 wire \dataBus[148] ;
 wire \dataBus[149] ;
 wire \dataBus[14] ;
 wire \dataBus[150] ;
 wire \dataBus[151] ;
 wire \dataBus[152] ;
 wire \dataBus[153] ;
 wire \dataBus[154] ;
 wire \dataBus[155] ;
 wire \dataBus[156] ;
 wire \dataBus[157] ;
 wire \dataBus[158] ;
 wire \dataBus[159] ;
 wire \dataBus[15] ;
 wire \dataBus[160] ;
 wire \dataBus[161] ;
 wire \dataBus[162] ;
 wire \dataBus[16] ;
 wire \dataBus[17] ;
 wire \dataBus[18] ;
 wire \dataBus[19] ;
 wire \dataBus[1] ;
 wire \dataBus[20] ;
 wire \dataBus[21] ;
 wire \dataBus[22] ;
 wire \dataBus[23] ;
 wire \dataBus[24] ;
 wire \dataBus[25] ;
 wire \dataBus[26] ;
 wire \dataBus[27] ;
 wire \dataBus[28] ;
 wire \dataBus[29] ;
 wire \dataBus[2] ;
 wire \dataBus[30] ;
 wire \dataBus[31] ;
 wire \dataBus[32] ;
 wire \dataBus[33] ;
 wire \dataBus[34] ;
 wire \dataBus[35] ;
 wire \dataBus[36] ;
 wire \dataBus[37] ;
 wire \dataBus[38] ;
 wire \dataBus[39] ;
 wire \dataBus[3] ;
 wire \dataBus[40] ;
 wire \dataBus[41] ;
 wire \dataBus[42] ;
 wire \dataBus[43] ;
 wire \dataBus[44] ;
 wire \dataBus[45] ;
 wire \dataBus[46] ;
 wire \dataBus[47] ;
 wire \dataBus[48] ;
 wire \dataBus[49] ;
 wire \dataBus[4] ;
 wire \dataBus[50] ;
 wire \dataBus[51] ;
 wire \dataBus[52] ;
 wire \dataBus[53] ;
 wire \dataBus[54] ;
 wire \dataBus[55] ;
 wire \dataBus[56] ;
 wire \dataBus[57] ;
 wire \dataBus[58] ;
 wire \dataBus[59] ;
 wire \dataBus[5] ;
 wire \dataBus[60] ;
 wire \dataBus[61] ;
 wire \dataBus[62] ;
 wire \dataBus[63] ;
 wire \dataBus[64] ;
 wire \dataBus[65] ;
 wire \dataBus[66] ;
 wire \dataBus[67] ;
 wire \dataBus[68] ;
 wire \dataBus[69] ;
 wire \dataBus[6] ;
 wire \dataBus[70] ;
 wire \dataBus[71] ;
 wire \dataBus[72] ;
 wire \dataBus[73] ;
 wire \dataBus[74] ;
 wire \dataBus[75] ;
 wire \dataBus[76] ;
 wire \dataBus[77] ;
 wire \dataBus[78] ;
 wire \dataBus[79] ;
 wire \dataBus[7] ;
 wire \dataBus[80] ;
 wire \dataBus[81] ;
 wire \dataBus[82] ;
 wire \dataBus[83] ;
 wire \dataBus[84] ;
 wire \dataBus[85] ;
 wire \dataBus[86] ;
 wire \dataBus[87] ;
 wire \dataBus[88] ;
 wire \dataBus[89] ;
 wire \dataBus[8] ;
 wire \dataBus[90] ;
 wire \dataBus[91] ;
 wire \dataBus[92] ;
 wire \dataBus[93] ;
 wire \dataBus[94] ;
 wire \dataBus[95] ;
 wire \dataBus[96] ;
 wire \dataBus[97] ;
 wire \dataBus[98] ;
 wire \dataBus[99] ;
 wire \dataBus[9] ;
 wire ki;
 wire next_key;
 wire slave_ena;
 wire \w_becStatus[0] ;
 wire \w_becStatus[1] ;
 wire \w_becStatus[2] ;
 wire \w_becStatus[3] ;
 wire \w_loadStatus[0] ;
 wire \w_loadStatus[1] ;
 wire \w_loadStatus[2] ;
 wire w_load_data;
 wire w_slvDone;
 wire w_trigLoad;

 sm_bec_v3 bec_core (.clk(wb_clk_i),
    .done(w_slvDone),
    .enable(slave_ena),
    .ki(ki),
    .load_data(w_load_data),
    .next_key(next_key),
    .rst(wb_rst_i),
    .trigLoad(w_trigLoad),
    .becStatus({\w_becStatus[3] ,
    \w_becStatus[2] ,
    \w_becStatus[1] ,
    \w_becStatus[0] }),
    .data_in({\configBus[162] ,
    \configBus[161] ,
    \configBus[160] ,
    \configBus[159] ,
    \configBus[158] ,
    \configBus[157] ,
    \configBus[156] ,
    \configBus[155] ,
    \configBus[154] ,
    \configBus[153] ,
    \configBus[152] ,
    \configBus[151] ,
    \configBus[150] ,
    \configBus[149] ,
    \configBus[148] ,
    \configBus[147] ,
    \configBus[146] ,
    \configBus[145] ,
    \configBus[144] ,
    \configBus[143] ,
    \configBus[142] ,
    \configBus[141] ,
    \configBus[140] ,
    \configBus[139] ,
    \configBus[138] ,
    \configBus[137] ,
    \configBus[136] ,
    \configBus[135] ,
    \configBus[134] ,
    \configBus[133] ,
    \configBus[132] ,
    \configBus[131] ,
    \configBus[130] ,
    \configBus[129] ,
    \configBus[128] ,
    \configBus[127] ,
    \configBus[126] ,
    \configBus[125] ,
    \configBus[124] ,
    \configBus[123] ,
    \configBus[122] ,
    \configBus[121] ,
    \configBus[120] ,
    \configBus[119] ,
    \configBus[118] ,
    \configBus[117] ,
    \configBus[116] ,
    \configBus[115] ,
    \configBus[114] ,
    \configBus[113] ,
    \configBus[112] ,
    \configBus[111] ,
    \configBus[110] ,
    \configBus[109] ,
    \configBus[108] ,
    \configBus[107] ,
    \configBus[106] ,
    \configBus[105] ,
    \configBus[104] ,
    \configBus[103] ,
    \configBus[102] ,
    \configBus[101] ,
    \configBus[100] ,
    \configBus[99] ,
    \configBus[98] ,
    \configBus[97] ,
    \configBus[96] ,
    \configBus[95] ,
    \configBus[94] ,
    \configBus[93] ,
    \configBus[92] ,
    \configBus[91] ,
    \configBus[90] ,
    \configBus[89] ,
    \configBus[88] ,
    \configBus[87] ,
    \configBus[86] ,
    \configBus[85] ,
    \configBus[84] ,
    \configBus[83] ,
    \configBus[82] ,
    \configBus[81] ,
    \configBus[80] ,
    \configBus[79] ,
    \configBus[78] ,
    \configBus[77] ,
    \configBus[76] ,
    \configBus[75] ,
    \configBus[74] ,
    \configBus[73] ,
    \configBus[72] ,
    \configBus[71] ,
    \configBus[70] ,
    \configBus[69] ,
    \configBus[68] ,
    \configBus[67] ,
    \configBus[66] ,
    \configBus[65] ,
    \configBus[64] ,
    \configBus[63] ,
    \configBus[62] ,
    \configBus[61] ,
    \configBus[60] ,
    \configBus[59] ,
    \configBus[58] ,
    \configBus[57] ,
    \configBus[56] ,
    \configBus[55] ,
    \configBus[54] ,
    \configBus[53] ,
    \configBus[52] ,
    \configBus[51] ,
    \configBus[50] ,
    \configBus[49] ,
    \configBus[48] ,
    \configBus[47] ,
    \configBus[46] ,
    \configBus[45] ,
    \configBus[44] ,
    \configBus[43] ,
    \configBus[42] ,
    \configBus[41] ,
    \configBus[40] ,
    \configBus[39] ,
    \configBus[38] ,
    \configBus[37] ,
    \configBus[36] ,
    \configBus[35] ,
    \configBus[34] ,
    \configBus[33] ,
    \configBus[32] ,
    \configBus[31] ,
    \configBus[30] ,
    \configBus[29] ,
    \configBus[28] ,
    \configBus[27] ,
    \configBus[26] ,
    \configBus[25] ,
    \configBus[24] ,
    \configBus[23] ,
    \configBus[22] ,
    \configBus[21] ,
    \configBus[20] ,
    \configBus[19] ,
    \configBus[18] ,
    \configBus[17] ,
    \configBus[16] ,
    \configBus[15] ,
    \configBus[14] ,
    \configBus[13] ,
    \configBus[12] ,
    \configBus[11] ,
    \configBus[10] ,
    \configBus[9] ,
    \configBus[8] ,
    \configBus[7] ,
    \configBus[6] ,
    \configBus[5] ,
    \configBus[4] ,
    \configBus[3] ,
    \configBus[2] ,
    \configBus[1] ,
    \configBus[0] }),
    .data_out({\dataBus[162] ,
    \dataBus[161] ,
    \dataBus[160] ,
    \dataBus[159] ,
    \dataBus[158] ,
    \dataBus[157] ,
    \dataBus[156] ,
    \dataBus[155] ,
    \dataBus[154] ,
    \dataBus[153] ,
    \dataBus[152] ,
    \dataBus[151] ,
    \dataBus[150] ,
    \dataBus[149] ,
    \dataBus[148] ,
    \dataBus[147] ,
    \dataBus[146] ,
    \dataBus[145] ,
    \dataBus[144] ,
    \dataBus[143] ,
    \dataBus[142] ,
    \dataBus[141] ,
    \dataBus[140] ,
    \dataBus[139] ,
    \dataBus[138] ,
    \dataBus[137] ,
    \dataBus[136] ,
    \dataBus[135] ,
    \dataBus[134] ,
    \dataBus[133] ,
    \dataBus[132] ,
    \dataBus[131] ,
    \dataBus[130] ,
    \dataBus[129] ,
    \dataBus[128] ,
    \dataBus[127] ,
    \dataBus[126] ,
    \dataBus[125] ,
    \dataBus[124] ,
    \dataBus[123] ,
    \dataBus[122] ,
    \dataBus[121] ,
    \dataBus[120] ,
    \dataBus[119] ,
    \dataBus[118] ,
    \dataBus[117] ,
    \dataBus[116] ,
    \dataBus[115] ,
    \dataBus[114] ,
    \dataBus[113] ,
    \dataBus[112] ,
    \dataBus[111] ,
    \dataBus[110] ,
    \dataBus[109] ,
    \dataBus[108] ,
    \dataBus[107] ,
    \dataBus[106] ,
    \dataBus[105] ,
    \dataBus[104] ,
    \dataBus[103] ,
    \dataBus[102] ,
    \dataBus[101] ,
    \dataBus[100] ,
    \dataBus[99] ,
    \dataBus[98] ,
    \dataBus[97] ,
    \dataBus[96] ,
    \dataBus[95] ,
    \dataBus[94] ,
    \dataBus[93] ,
    \dataBus[92] ,
    \dataBus[91] ,
    \dataBus[90] ,
    \dataBus[89] ,
    \dataBus[88] ,
    \dataBus[87] ,
    \dataBus[86] ,
    \dataBus[85] ,
    \dataBus[84] ,
    \dataBus[83] ,
    \dataBus[82] ,
    \dataBus[81] ,
    \dataBus[80] ,
    \dataBus[79] ,
    \dataBus[78] ,
    \dataBus[77] ,
    \dataBus[76] ,
    \dataBus[75] ,
    \dataBus[74] ,
    \dataBus[73] ,
    \dataBus[72] ,
    \dataBus[71] ,
    \dataBus[70] ,
    \dataBus[69] ,
    \dataBus[68] ,
    \dataBus[67] ,
    \dataBus[66] ,
    \dataBus[65] ,
    \dataBus[64] ,
    \dataBus[63] ,
    \dataBus[62] ,
    \dataBus[61] ,
    \dataBus[60] ,
    \dataBus[59] ,
    \dataBus[58] ,
    \dataBus[57] ,
    \dataBus[56] ,
    \dataBus[55] ,
    \dataBus[54] ,
    \dataBus[53] ,
    \dataBus[52] ,
    \dataBus[51] ,
    \dataBus[50] ,
    \dataBus[49] ,
    \dataBus[48] ,
    \dataBus[47] ,
    \dataBus[46] ,
    \dataBus[45] ,
    \dataBus[44] ,
    \dataBus[43] ,
    \dataBus[42] ,
    \dataBus[41] ,
    \dataBus[40] ,
    \dataBus[39] ,
    \dataBus[38] ,
    \dataBus[37] ,
    \dataBus[36] ,
    \dataBus[35] ,
    \dataBus[34] ,
    \dataBus[33] ,
    \dataBus[32] ,
    \dataBus[31] ,
    \dataBus[30] ,
    \dataBus[29] ,
    \dataBus[28] ,
    \dataBus[27] ,
    \dataBus[26] ,
    \dataBus[25] ,
    \dataBus[24] ,
    \dataBus[23] ,
    \dataBus[22] ,
    \dataBus[21] ,
    \dataBus[20] ,
    \dataBus[19] ,
    \dataBus[18] ,
    \dataBus[17] ,
    \dataBus[16] ,
    \dataBus[15] ,
    \dataBus[14] ,
    \dataBus[13] ,
    \dataBus[12] ,
    \dataBus[11] ,
    \dataBus[10] ,
    \dataBus[9] ,
    \dataBus[8] ,
    \dataBus[7] ,
    \dataBus[6] ,
    \dataBus[5] ,
    \dataBus[4] ,
    \dataBus[3] ,
    \dataBus[2] ,
    \dataBus[1] ,
    \dataBus[0] }),
    .load_status({\w_loadStatus[2] ,
    \w_loadStatus[1] ,
    \w_loadStatus[0] }));
 controller control_unit (.ki(ki),
    .load_data(w_load_data),
    .master_ena_proc(slave_ena),
    .next_key(next_key),
    .slv_done(w_slvDone),
    .trigLoad(w_trigLoad),
    .wb_clk_i(wb_clk_i),
    .wb_rst_i(wb_rst_i),
    .becStatus({\w_becStatus[3] ,
    \w_becStatus[2] ,
    \w_becStatus[1] ,
    \w_becStatus[0] }),
    .data_in({\dataBus[162] ,
    \dataBus[161] ,
    \dataBus[160] ,
    \dataBus[159] ,
    \dataBus[158] ,
    \dataBus[157] ,
    \dataBus[156] ,
    \dataBus[155] ,
    \dataBus[154] ,
    \dataBus[153] ,
    \dataBus[152] ,
    \dataBus[151] ,
    \dataBus[150] ,
    \dataBus[149] ,
    \dataBus[148] ,
    \dataBus[147] ,
    \dataBus[146] ,
    \dataBus[145] ,
    \dataBus[144] ,
    \dataBus[143] ,
    \dataBus[142] ,
    \dataBus[141] ,
    \dataBus[140] ,
    \dataBus[139] ,
    \dataBus[138] ,
    \dataBus[137] ,
    \dataBus[136] ,
    \dataBus[135] ,
    \dataBus[134] ,
    \dataBus[133] ,
    \dataBus[132] ,
    \dataBus[131] ,
    \dataBus[130] ,
    \dataBus[129] ,
    \dataBus[128] ,
    \dataBus[127] ,
    \dataBus[126] ,
    \dataBus[125] ,
    \dataBus[124] ,
    \dataBus[123] ,
    \dataBus[122] ,
    \dataBus[121] ,
    \dataBus[120] ,
    \dataBus[119] ,
    \dataBus[118] ,
    \dataBus[117] ,
    \dataBus[116] ,
    \dataBus[115] ,
    \dataBus[114] ,
    \dataBus[113] ,
    \dataBus[112] ,
    \dataBus[111] ,
    \dataBus[110] ,
    \dataBus[109] ,
    \dataBus[108] ,
    \dataBus[107] ,
    \dataBus[106] ,
    \dataBus[105] ,
    \dataBus[104] ,
    \dataBus[103] ,
    \dataBus[102] ,
    \dataBus[101] ,
    \dataBus[100] ,
    \dataBus[99] ,
    \dataBus[98] ,
    \dataBus[97] ,
    \dataBus[96] ,
    \dataBus[95] ,
    \dataBus[94] ,
    \dataBus[93] ,
    \dataBus[92] ,
    \dataBus[91] ,
    \dataBus[90] ,
    \dataBus[89] ,
    \dataBus[88] ,
    \dataBus[87] ,
    \dataBus[86] ,
    \dataBus[85] ,
    \dataBus[84] ,
    \dataBus[83] ,
    \dataBus[82] ,
    \dataBus[81] ,
    \dataBus[80] ,
    \dataBus[79] ,
    \dataBus[78] ,
    \dataBus[77] ,
    \dataBus[76] ,
    \dataBus[75] ,
    \dataBus[74] ,
    \dataBus[73] ,
    \dataBus[72] ,
    \dataBus[71] ,
    \dataBus[70] ,
    \dataBus[69] ,
    \dataBus[68] ,
    \dataBus[67] ,
    \dataBus[66] ,
    \dataBus[65] ,
    \dataBus[64] ,
    \dataBus[63] ,
    \dataBus[62] ,
    \dataBus[61] ,
    \dataBus[60] ,
    \dataBus[59] ,
    \dataBus[58] ,
    \dataBus[57] ,
    \dataBus[56] ,
    \dataBus[55] ,
    \dataBus[54] ,
    \dataBus[53] ,
    \dataBus[52] ,
    \dataBus[51] ,
    \dataBus[50] ,
    \dataBus[49] ,
    \dataBus[48] ,
    \dataBus[47] ,
    \dataBus[46] ,
    \dataBus[45] ,
    \dataBus[44] ,
    \dataBus[43] ,
    \dataBus[42] ,
    \dataBus[41] ,
    \dataBus[40] ,
    \dataBus[39] ,
    \dataBus[38] ,
    \dataBus[37] ,
    \dataBus[36] ,
    \dataBus[35] ,
    \dataBus[34] ,
    \dataBus[33] ,
    \dataBus[32] ,
    \dataBus[31] ,
    \dataBus[30] ,
    \dataBus[29] ,
    \dataBus[28] ,
    \dataBus[27] ,
    \dataBus[26] ,
    \dataBus[25] ,
    \dataBus[24] ,
    \dataBus[23] ,
    \dataBus[22] ,
    \dataBus[21] ,
    \dataBus[20] ,
    \dataBus[19] ,
    \dataBus[18] ,
    \dataBus[17] ,
    \dataBus[16] ,
    \dataBus[15] ,
    \dataBus[14] ,
    \dataBus[13] ,
    \dataBus[12] ,
    \dataBus[11] ,
    \dataBus[10] ,
    \dataBus[9] ,
    \dataBus[8] ,
    \dataBus[7] ,
    \dataBus[6] ,
    \dataBus[5] ,
    \dataBus[4] ,
    \dataBus[3] ,
    \dataBus[2] ,
    \dataBus[1] ,
    \dataBus[0] }),
    .data_out({\configBus[162] ,
    \configBus[161] ,
    \configBus[160] ,
    \configBus[159] ,
    \configBus[158] ,
    \configBus[157] ,
    \configBus[156] ,
    \configBus[155] ,
    \configBus[154] ,
    \configBus[153] ,
    \configBus[152] ,
    \configBus[151] ,
    \configBus[150] ,
    \configBus[149] ,
    \configBus[148] ,
    \configBus[147] ,
    \configBus[146] ,
    \configBus[145] ,
    \configBus[144] ,
    \configBus[143] ,
    \configBus[142] ,
    \configBus[141] ,
    \configBus[140] ,
    \configBus[139] ,
    \configBus[138] ,
    \configBus[137] ,
    \configBus[136] ,
    \configBus[135] ,
    \configBus[134] ,
    \configBus[133] ,
    \configBus[132] ,
    \configBus[131] ,
    \configBus[130] ,
    \configBus[129] ,
    \configBus[128] ,
    \configBus[127] ,
    \configBus[126] ,
    \configBus[125] ,
    \configBus[124] ,
    \configBus[123] ,
    \configBus[122] ,
    \configBus[121] ,
    \configBus[120] ,
    \configBus[119] ,
    \configBus[118] ,
    \configBus[117] ,
    \configBus[116] ,
    \configBus[115] ,
    \configBus[114] ,
    \configBus[113] ,
    \configBus[112] ,
    \configBus[111] ,
    \configBus[110] ,
    \configBus[109] ,
    \configBus[108] ,
    \configBus[107] ,
    \configBus[106] ,
    \configBus[105] ,
    \configBus[104] ,
    \configBus[103] ,
    \configBus[102] ,
    \configBus[101] ,
    \configBus[100] ,
    \configBus[99] ,
    \configBus[98] ,
    \configBus[97] ,
    \configBus[96] ,
    \configBus[95] ,
    \configBus[94] ,
    \configBus[93] ,
    \configBus[92] ,
    \configBus[91] ,
    \configBus[90] ,
    \configBus[89] ,
    \configBus[88] ,
    \configBus[87] ,
    \configBus[86] ,
    \configBus[85] ,
    \configBus[84] ,
    \configBus[83] ,
    \configBus[82] ,
    \configBus[81] ,
    \configBus[80] ,
    \configBus[79] ,
    \configBus[78] ,
    \configBus[77] ,
    \configBus[76] ,
    \configBus[75] ,
    \configBus[74] ,
    \configBus[73] ,
    \configBus[72] ,
    \configBus[71] ,
    \configBus[70] ,
    \configBus[69] ,
    \configBus[68] ,
    \configBus[67] ,
    \configBus[66] ,
    \configBus[65] ,
    \configBus[64] ,
    \configBus[63] ,
    \configBus[62] ,
    \configBus[61] ,
    \configBus[60] ,
    \configBus[59] ,
    \configBus[58] ,
    \configBus[57] ,
    \configBus[56] ,
    \configBus[55] ,
    \configBus[54] ,
    \configBus[53] ,
    \configBus[52] ,
    \configBus[51] ,
    \configBus[50] ,
    \configBus[49] ,
    \configBus[48] ,
    \configBus[47] ,
    \configBus[46] ,
    \configBus[45] ,
    \configBus[44] ,
    \configBus[43] ,
    \configBus[42] ,
    \configBus[41] ,
    \configBus[40] ,
    \configBus[39] ,
    \configBus[38] ,
    \configBus[37] ,
    \configBus[36] ,
    \configBus[35] ,
    \configBus[34] ,
    \configBus[33] ,
    \configBus[32] ,
    \configBus[31] ,
    \configBus[30] ,
    \configBus[29] ,
    \configBus[28] ,
    \configBus[27] ,
    \configBus[26] ,
    \configBus[25] ,
    \configBus[24] ,
    \configBus[23] ,
    \configBus[22] ,
    \configBus[21] ,
    \configBus[20] ,
    \configBus[19] ,
    \configBus[18] ,
    \configBus[17] ,
    \configBus[16] ,
    \configBus[15] ,
    \configBus[14] ,
    \configBus[13] ,
    \configBus[12] ,
    \configBus[11] ,
    \configBus[10] ,
    \configBus[9] ,
    \configBus[8] ,
    \configBus[7] ,
    \configBus[6] ,
    \configBus[5] ,
    \configBus[4] ,
    \configBus[3] ,
    \configBus[2] ,
    \configBus[1] ,
    \configBus[0] }),
    .la_data_in({la_data_in[127],
    la_data_in[126],
    la_data_in[125],
    la_data_in[124],
    la_data_in[123],
    la_data_in[122],
    la_data_in[121],
    la_data_in[120],
    la_data_in[119],
    la_data_in[118],
    la_data_in[117],
    la_data_in[116],
    la_data_in[115],
    la_data_in[114],
    la_data_in[113],
    la_data_in[112],
    la_data_in[111],
    la_data_in[110],
    la_data_in[109],
    la_data_in[108],
    la_data_in[107],
    la_data_in[106],
    la_data_in[105],
    la_data_in[104],
    la_data_in[103],
    la_data_in[102],
    la_data_in[101],
    la_data_in[100],
    la_data_in[99],
    la_data_in[98],
    la_data_in[97],
    la_data_in[96],
    la_data_in[95],
    la_data_in[94],
    la_data_in[93],
    la_data_in[92],
    la_data_in[91],
    la_data_in[90],
    la_data_in[89],
    la_data_in[88],
    la_data_in[87],
    la_data_in[86],
    la_data_in[85],
    la_data_in[84],
    la_data_in[83],
    la_data_in[82],
    la_data_in[81],
    la_data_in[80],
    la_data_in[79],
    la_data_in[78],
    la_data_in[77],
    la_data_in[76],
    la_data_in[75],
    la_data_in[74],
    la_data_in[73],
    la_data_in[72],
    la_data_in[71],
    la_data_in[70],
    la_data_in[69],
    la_data_in[68],
    la_data_in[67],
    la_data_in[66],
    la_data_in[65],
    la_data_in[64],
    la_data_in[63],
    la_data_in[62],
    la_data_in[61],
    la_data_in[60],
    la_data_in[59],
    la_data_in[58],
    la_data_in[57],
    la_data_in[56],
    la_data_in[55],
    la_data_in[54],
    la_data_in[53],
    la_data_in[52],
    la_data_in[51],
    la_data_in[50],
    la_data_in[49],
    la_data_in[48],
    la_data_in[47],
    la_data_in[46],
    la_data_in[45],
    la_data_in[44],
    la_data_in[43],
    la_data_in[42],
    la_data_in[41],
    la_data_in[40],
    la_data_in[39],
    la_data_in[38],
    la_data_in[37],
    la_data_in[36],
    la_data_in[35],
    la_data_in[34],
    la_data_in[33],
    la_data_in[32],
    la_data_in[31],
    la_data_in[30],
    la_data_in[29],
    la_data_in[28],
    la_data_in[27],
    la_data_in[26],
    la_data_in[25],
    la_data_in[24],
    la_data_in[23],
    la_data_in[22],
    la_data_in[21],
    la_data_in[20],
    la_data_in[19],
    la_data_in[18],
    la_data_in[17],
    la_data_in[16],
    la_data_in[15],
    la_data_in[14],
    la_data_in[13],
    la_data_in[12],
    la_data_in[11],
    la_data_in[10],
    la_data_in[9],
    la_data_in[8],
    la_data_in[7],
    la_data_in[6],
    la_data_in[5],
    la_data_in[4],
    la_data_in[3],
    la_data_in[2],
    la_data_in[1],
    la_data_in[0]}),
    .la_data_out({la_data_out[127],
    la_data_out[126],
    la_data_out[125],
    la_data_out[124],
    la_data_out[123],
    la_data_out[122],
    la_data_out[121],
    la_data_out[120],
    la_data_out[119],
    la_data_out[118],
    la_data_out[117],
    la_data_out[116],
    la_data_out[115],
    la_data_out[114],
    la_data_out[113],
    la_data_out[112],
    la_data_out[111],
    la_data_out[110],
    la_data_out[109],
    la_data_out[108],
    la_data_out[107],
    la_data_out[106],
    la_data_out[105],
    la_data_out[104],
    la_data_out[103],
    la_data_out[102],
    la_data_out[101],
    la_data_out[100],
    la_data_out[99],
    la_data_out[98],
    la_data_out[97],
    la_data_out[96],
    la_data_out[95],
    la_data_out[94],
    la_data_out[93],
    la_data_out[92],
    la_data_out[91],
    la_data_out[90],
    la_data_out[89],
    la_data_out[88],
    la_data_out[87],
    la_data_out[86],
    la_data_out[85],
    la_data_out[84],
    la_data_out[83],
    la_data_out[82],
    la_data_out[81],
    la_data_out[80],
    la_data_out[79],
    la_data_out[78],
    la_data_out[77],
    la_data_out[76],
    la_data_out[75],
    la_data_out[74],
    la_data_out[73],
    la_data_out[72],
    la_data_out[71],
    la_data_out[70],
    la_data_out[69],
    la_data_out[68],
    la_data_out[67],
    la_data_out[66],
    la_data_out[65],
    la_data_out[64],
    la_data_out[63],
    la_data_out[62],
    la_data_out[61],
    la_data_out[60],
    la_data_out[59],
    la_data_out[58],
    la_data_out[57],
    la_data_out[56],
    la_data_out[55],
    la_data_out[54],
    la_data_out[53],
    la_data_out[52],
    la_data_out[51],
    la_data_out[50],
    la_data_out[49],
    la_data_out[48],
    la_data_out[47],
    la_data_out[46],
    la_data_out[45],
    la_data_out[44],
    la_data_out[43],
    la_data_out[42],
    la_data_out[41],
    la_data_out[40],
    la_data_out[39],
    la_data_out[38],
    la_data_out[37],
    la_data_out[36],
    la_data_out[35],
    la_data_out[34],
    la_data_out[33],
    la_data_out[32],
    la_data_out[31],
    la_data_out[30],
    la_data_out[29],
    la_data_out[28],
    la_data_out[27],
    la_data_out[26],
    la_data_out[25],
    la_data_out[24],
    la_data_out[23],
    la_data_out[22],
    la_data_out[21],
    la_data_out[20],
    la_data_out[19],
    la_data_out[18],
    la_data_out[17],
    la_data_out[16],
    la_data_out[15],
    la_data_out[14],
    la_data_out[13],
    la_data_out[12],
    la_data_out[11],
    la_data_out[10],
    la_data_out[9],
    la_data_out[8],
    la_data_out[7],
    la_data_out[6],
    la_data_out[5],
    la_data_out[4],
    la_data_out[3],
    la_data_out[2],
    la_data_out[1],
    la_data_out[0]}),
    .la_oenb({la_oenb[127],
    la_oenb[126],
    la_oenb[125],
    la_oenb[124],
    la_oenb[123],
    la_oenb[122],
    la_oenb[121],
    la_oenb[120],
    la_oenb[119],
    la_oenb[118],
    la_oenb[117],
    la_oenb[116],
    la_oenb[115],
    la_oenb[114],
    la_oenb[113],
    la_oenb[112],
    la_oenb[111],
    la_oenb[110],
    la_oenb[109],
    la_oenb[108],
    la_oenb[107],
    la_oenb[106],
    la_oenb[105],
    la_oenb[104],
    la_oenb[103],
    la_oenb[102],
    la_oenb[101],
    la_oenb[100],
    la_oenb[99],
    la_oenb[98],
    la_oenb[97],
    la_oenb[96],
    la_oenb[95],
    la_oenb[94],
    la_oenb[93],
    la_oenb[92],
    la_oenb[91],
    la_oenb[90],
    la_oenb[89],
    la_oenb[88],
    la_oenb[87],
    la_oenb[86],
    la_oenb[85],
    la_oenb[84],
    la_oenb[83],
    la_oenb[82],
    la_oenb[81],
    la_oenb[80],
    la_oenb[79],
    la_oenb[78],
    la_oenb[77],
    la_oenb[76],
    la_oenb[75],
    la_oenb[74],
    la_oenb[73],
    la_oenb[72],
    la_oenb[71],
    la_oenb[70],
    la_oenb[69],
    la_oenb[68],
    la_oenb[67],
    la_oenb[66],
    la_oenb[65],
    la_oenb[64],
    la_oenb[63],
    la_oenb[62],
    la_oenb[61],
    la_oenb[60],
    la_oenb[59],
    la_oenb[58],
    la_oenb[57],
    la_oenb[56],
    la_oenb[55],
    la_oenb[54],
    la_oenb[53],
    la_oenb[52],
    la_oenb[51],
    la_oenb[50],
    la_oenb[49],
    la_oenb[48],
    la_oenb[47],
    la_oenb[46],
    la_oenb[45],
    la_oenb[44],
    la_oenb[43],
    la_oenb[42],
    la_oenb[41],
    la_oenb[40],
    la_oenb[39],
    la_oenb[38],
    la_oenb[37],
    la_oenb[36],
    la_oenb[35],
    la_oenb[34],
    la_oenb[33],
    la_oenb[32],
    la_oenb[31],
    la_oenb[30],
    la_oenb[29],
    la_oenb[28],
    la_oenb[27],
    la_oenb[26],
    la_oenb[25],
    la_oenb[24],
    la_oenb[23],
    la_oenb[22],
    la_oenb[21],
    la_oenb[20],
    la_oenb[19],
    la_oenb[18],
    la_oenb[17],
    la_oenb[16],
    la_oenb[15],
    la_oenb[14],
    la_oenb[13],
    la_oenb[12],
    la_oenb[11],
    la_oenb[10],
    la_oenb[9],
    la_oenb[8],
    la_oenb[7],
    la_oenb[6],
    la_oenb[5],
    la_oenb[4],
    la_oenb[3],
    la_oenb[2],
    la_oenb[1],
    la_oenb[0]}),
    .load_status({\w_loadStatus[2] ,
    \w_loadStatus[1] ,
    \w_loadStatus[0] }));
endmodule

