// SPDX-FileCopyrightText: 2020 Efabless Corporation
//
// Licensed under the Apache License, Version 2.0 (the "License");
// you may not use this file except in compliance with the License.
// You may obtain a copy of the License at
//
//      http://www.apache.org/licenses/LICENSE-2.0
//
// Unless required by applicable law or agreed to in writing, software
// distributed under the License is distributed on an "AS IS" BASIS,
// WITHOUT WARRANTIES OR CONDITIONS OF ANY KIND, either express or implied.
// See the License for the specific language governing permissions and
// limitations under the License.
// SPDX-License-Identifier: Apache-2.0

// `default_nettype none
//`include "../../../verilog/rtl/classic_squarer.v"
//`include "../../../verilog/rtl/interleaved_mult.v"

module acb (
    `ifdef USE_POWER_PINS
        inout vccd2,	// User area 2 1.8v supply
        inout vssd2,	// User area 2 digital ground
    `endif
    
    clk, rst, enable, configuration, A, B, C, done);
    input clk, rst, enable, configuration;
    input [162:0] A, B;

    output wire [162:0] C;

    output wire done;

    wire [162:0] z_tmp, c_tmp;
    assign C = (~configuration) ? c_tmp : z_tmp; 

    classic_squarer u1 (
        .a(z_tmp),
        .c(c_tmp)
    );

    interleaved_mult u2 (
        `ifdef USE_POWER_PINS
			.vccd2(vccd2),	// User area 2 1.8v supply
			.vssd2(vssd2),	// User area 2 digital ground
		`endif
        .A(A),
        .B(B),
        .clk(clk),
        .rst(rst),
        .start(enable),
        .Z(z_tmp),
        .done(done)
    );

    // always @(posedge clk or rst) begin
    //     if (rst) begin
    //         C <= 0;
    //     end else begin
    //         if (~configuration)
    //             C <= c_tmp;
    //         else
    //             C <= z_tmp;
    //     end
    // end
endmodule
`default_nettype wire
